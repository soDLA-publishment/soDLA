module NV_NVDLA_CMAC_CORE_rt_in(
  input        clock,
  input        reset,
  input  [7:0] io_sc2mac_dat_data_0,
  input  [7:0] io_sc2mac_dat_data_1,
  input  [7:0] io_sc2mac_dat_data_2,
  input  [7:0] io_sc2mac_dat_data_3,
  input  [7:0] io_sc2mac_dat_data_4,
  input  [7:0] io_sc2mac_dat_data_5,
  input  [7:0] io_sc2mac_dat_data_6,
  input  [7:0] io_sc2mac_dat_data_7,
  input  [7:0] io_sc2mac_dat_data_8,
  input  [7:0] io_sc2mac_dat_data_9,
  input  [7:0] io_sc2mac_dat_data_10,
  input  [7:0] io_sc2mac_dat_data_11,
  input  [7:0] io_sc2mac_dat_data_12,
  input  [7:0] io_sc2mac_dat_data_13,
  input  [7:0] io_sc2mac_dat_data_14,
  input  [7:0] io_sc2mac_dat_data_15,
  input  [7:0] io_sc2mac_dat_data_16,
  input  [7:0] io_sc2mac_dat_data_17,
  input  [7:0] io_sc2mac_dat_data_18,
  input  [7:0] io_sc2mac_dat_data_19,
  input  [7:0] io_sc2mac_dat_data_20,
  input  [7:0] io_sc2mac_dat_data_21,
  input  [7:0] io_sc2mac_dat_data_22,
  input  [7:0] io_sc2mac_dat_data_23,
  input  [7:0] io_sc2mac_dat_data_24,
  input  [7:0] io_sc2mac_dat_data_25,
  input  [7:0] io_sc2mac_dat_data_26,
  input  [7:0] io_sc2mac_dat_data_27,
  input  [7:0] io_sc2mac_dat_data_28,
  input  [7:0] io_sc2mac_dat_data_29,
  input  [7:0] io_sc2mac_dat_data_30,
  input  [7:0] io_sc2mac_dat_data_31,
  input  [7:0] io_sc2mac_dat_data_32,
  input  [7:0] io_sc2mac_dat_data_33,
  input  [7:0] io_sc2mac_dat_data_34,
  input  [7:0] io_sc2mac_dat_data_35,
  input  [7:0] io_sc2mac_dat_data_36,
  input  [7:0] io_sc2mac_dat_data_37,
  input  [7:0] io_sc2mac_dat_data_38,
  input  [7:0] io_sc2mac_dat_data_39,
  input  [7:0] io_sc2mac_dat_data_40,
  input  [7:0] io_sc2mac_dat_data_41,
  input  [7:0] io_sc2mac_dat_data_42,
  input  [7:0] io_sc2mac_dat_data_43,
  input  [7:0] io_sc2mac_dat_data_44,
  input  [7:0] io_sc2mac_dat_data_45,
  input  [7:0] io_sc2mac_dat_data_46,
  input  [7:0] io_sc2mac_dat_data_47,
  input  [7:0] io_sc2mac_dat_data_48,
  input  [7:0] io_sc2mac_dat_data_49,
  input  [7:0] io_sc2mac_dat_data_50,
  input  [7:0] io_sc2mac_dat_data_51,
  input  [7:0] io_sc2mac_dat_data_52,
  input  [7:0] io_sc2mac_dat_data_53,
  input  [7:0] io_sc2mac_dat_data_54,
  input  [7:0] io_sc2mac_dat_data_55,
  input  [7:0] io_sc2mac_dat_data_56,
  input  [7:0] io_sc2mac_dat_data_57,
  input  [7:0] io_sc2mac_dat_data_58,
  input  [7:0] io_sc2mac_dat_data_59,
  input  [7:0] io_sc2mac_dat_data_60,
  input  [7:0] io_sc2mac_dat_data_61,
  input  [7:0] io_sc2mac_dat_data_62,
  input  [7:0] io_sc2mac_dat_data_63,
  input  [7:0] io_sc2mac_dat_data_64,
  input  [7:0] io_sc2mac_dat_data_65,
  input  [7:0] io_sc2mac_dat_data_66,
  input  [7:0] io_sc2mac_dat_data_67,
  input  [7:0] io_sc2mac_dat_data_68,
  input  [7:0] io_sc2mac_dat_data_69,
  input  [7:0] io_sc2mac_dat_data_70,
  input  [7:0] io_sc2mac_dat_data_71,
  input  [7:0] io_sc2mac_dat_data_72,
  input  [7:0] io_sc2mac_dat_data_73,
  input  [7:0] io_sc2mac_dat_data_74,
  input  [7:0] io_sc2mac_dat_data_75,
  input  [7:0] io_sc2mac_dat_data_76,
  input  [7:0] io_sc2mac_dat_data_77,
  input  [7:0] io_sc2mac_dat_data_78,
  input  [7:0] io_sc2mac_dat_data_79,
  input  [7:0] io_sc2mac_dat_data_80,
  input  [7:0] io_sc2mac_dat_data_81,
  input  [7:0] io_sc2mac_dat_data_82,
  input  [7:0] io_sc2mac_dat_data_83,
  input  [7:0] io_sc2mac_dat_data_84,
  input  [7:0] io_sc2mac_dat_data_85,
  input  [7:0] io_sc2mac_dat_data_86,
  input  [7:0] io_sc2mac_dat_data_87,
  input  [7:0] io_sc2mac_dat_data_88,
  input  [7:0] io_sc2mac_dat_data_89,
  input  [7:0] io_sc2mac_dat_data_90,
  input  [7:0] io_sc2mac_dat_data_91,
  input  [7:0] io_sc2mac_dat_data_92,
  input  [7:0] io_sc2mac_dat_data_93,
  input  [7:0] io_sc2mac_dat_data_94,
  input  [7:0] io_sc2mac_dat_data_95,
  input  [7:0] io_sc2mac_dat_data_96,
  input  [7:0] io_sc2mac_dat_data_97,
  input  [7:0] io_sc2mac_dat_data_98,
  input  [7:0] io_sc2mac_dat_data_99,
  input  [7:0] io_sc2mac_dat_data_100,
  input  [7:0] io_sc2mac_dat_data_101,
  input  [7:0] io_sc2mac_dat_data_102,
  input  [7:0] io_sc2mac_dat_data_103,
  input  [7:0] io_sc2mac_dat_data_104,
  input  [7:0] io_sc2mac_dat_data_105,
  input  [7:0] io_sc2mac_dat_data_106,
  input  [7:0] io_sc2mac_dat_data_107,
  input  [7:0] io_sc2mac_dat_data_108,
  input  [7:0] io_sc2mac_dat_data_109,
  input  [7:0] io_sc2mac_dat_data_110,
  input  [7:0] io_sc2mac_dat_data_111,
  input  [7:0] io_sc2mac_dat_data_112,
  input  [7:0] io_sc2mac_dat_data_113,
  input  [7:0] io_sc2mac_dat_data_114,
  input  [7:0] io_sc2mac_dat_data_115,
  input  [7:0] io_sc2mac_dat_data_116,
  input  [7:0] io_sc2mac_dat_data_117,
  input  [7:0] io_sc2mac_dat_data_118,
  input  [7:0] io_sc2mac_dat_data_119,
  input  [7:0] io_sc2mac_dat_data_120,
  input  [7:0] io_sc2mac_dat_data_121,
  input  [7:0] io_sc2mac_dat_data_122,
  input  [7:0] io_sc2mac_dat_data_123,
  input  [7:0] io_sc2mac_dat_data_124,
  input  [7:0] io_sc2mac_dat_data_125,
  input  [7:0] io_sc2mac_dat_data_126,
  input  [7:0] io_sc2mac_dat_data_127,
  input        io_sc2mac_dat_mask_0,
  input        io_sc2mac_dat_mask_1,
  input        io_sc2mac_dat_mask_2,
  input        io_sc2mac_dat_mask_3,
  input        io_sc2mac_dat_mask_4,
  input        io_sc2mac_dat_mask_5,
  input        io_sc2mac_dat_mask_6,
  input        io_sc2mac_dat_mask_7,
  input        io_sc2mac_dat_mask_8,
  input        io_sc2mac_dat_mask_9,
  input        io_sc2mac_dat_mask_10,
  input        io_sc2mac_dat_mask_11,
  input        io_sc2mac_dat_mask_12,
  input        io_sc2mac_dat_mask_13,
  input        io_sc2mac_dat_mask_14,
  input        io_sc2mac_dat_mask_15,
  input        io_sc2mac_dat_mask_16,
  input        io_sc2mac_dat_mask_17,
  input        io_sc2mac_dat_mask_18,
  input        io_sc2mac_dat_mask_19,
  input        io_sc2mac_dat_mask_20,
  input        io_sc2mac_dat_mask_21,
  input        io_sc2mac_dat_mask_22,
  input        io_sc2mac_dat_mask_23,
  input        io_sc2mac_dat_mask_24,
  input        io_sc2mac_dat_mask_25,
  input        io_sc2mac_dat_mask_26,
  input        io_sc2mac_dat_mask_27,
  input        io_sc2mac_dat_mask_28,
  input        io_sc2mac_dat_mask_29,
  input        io_sc2mac_dat_mask_30,
  input        io_sc2mac_dat_mask_31,
  input        io_sc2mac_dat_mask_32,
  input        io_sc2mac_dat_mask_33,
  input        io_sc2mac_dat_mask_34,
  input        io_sc2mac_dat_mask_35,
  input        io_sc2mac_dat_mask_36,
  input        io_sc2mac_dat_mask_37,
  input        io_sc2mac_dat_mask_38,
  input        io_sc2mac_dat_mask_39,
  input        io_sc2mac_dat_mask_40,
  input        io_sc2mac_dat_mask_41,
  input        io_sc2mac_dat_mask_42,
  input        io_sc2mac_dat_mask_43,
  input        io_sc2mac_dat_mask_44,
  input        io_sc2mac_dat_mask_45,
  input        io_sc2mac_dat_mask_46,
  input        io_sc2mac_dat_mask_47,
  input        io_sc2mac_dat_mask_48,
  input        io_sc2mac_dat_mask_49,
  input        io_sc2mac_dat_mask_50,
  input        io_sc2mac_dat_mask_51,
  input        io_sc2mac_dat_mask_52,
  input        io_sc2mac_dat_mask_53,
  input        io_sc2mac_dat_mask_54,
  input        io_sc2mac_dat_mask_55,
  input        io_sc2mac_dat_mask_56,
  input        io_sc2mac_dat_mask_57,
  input        io_sc2mac_dat_mask_58,
  input        io_sc2mac_dat_mask_59,
  input        io_sc2mac_dat_mask_60,
  input        io_sc2mac_dat_mask_61,
  input        io_sc2mac_dat_mask_62,
  input        io_sc2mac_dat_mask_63,
  input        io_sc2mac_dat_mask_64,
  input        io_sc2mac_dat_mask_65,
  input        io_sc2mac_dat_mask_66,
  input        io_sc2mac_dat_mask_67,
  input        io_sc2mac_dat_mask_68,
  input        io_sc2mac_dat_mask_69,
  input        io_sc2mac_dat_mask_70,
  input        io_sc2mac_dat_mask_71,
  input        io_sc2mac_dat_mask_72,
  input        io_sc2mac_dat_mask_73,
  input        io_sc2mac_dat_mask_74,
  input        io_sc2mac_dat_mask_75,
  input        io_sc2mac_dat_mask_76,
  input        io_sc2mac_dat_mask_77,
  input        io_sc2mac_dat_mask_78,
  input        io_sc2mac_dat_mask_79,
  input        io_sc2mac_dat_mask_80,
  input        io_sc2mac_dat_mask_81,
  input        io_sc2mac_dat_mask_82,
  input        io_sc2mac_dat_mask_83,
  input        io_sc2mac_dat_mask_84,
  input        io_sc2mac_dat_mask_85,
  input        io_sc2mac_dat_mask_86,
  input        io_sc2mac_dat_mask_87,
  input        io_sc2mac_dat_mask_88,
  input        io_sc2mac_dat_mask_89,
  input        io_sc2mac_dat_mask_90,
  input        io_sc2mac_dat_mask_91,
  input        io_sc2mac_dat_mask_92,
  input        io_sc2mac_dat_mask_93,
  input        io_sc2mac_dat_mask_94,
  input        io_sc2mac_dat_mask_95,
  input        io_sc2mac_dat_mask_96,
  input        io_sc2mac_dat_mask_97,
  input        io_sc2mac_dat_mask_98,
  input        io_sc2mac_dat_mask_99,
  input        io_sc2mac_dat_mask_100,
  input        io_sc2mac_dat_mask_101,
  input        io_sc2mac_dat_mask_102,
  input        io_sc2mac_dat_mask_103,
  input        io_sc2mac_dat_mask_104,
  input        io_sc2mac_dat_mask_105,
  input        io_sc2mac_dat_mask_106,
  input        io_sc2mac_dat_mask_107,
  input        io_sc2mac_dat_mask_108,
  input        io_sc2mac_dat_mask_109,
  input        io_sc2mac_dat_mask_110,
  input        io_sc2mac_dat_mask_111,
  input        io_sc2mac_dat_mask_112,
  input        io_sc2mac_dat_mask_113,
  input        io_sc2mac_dat_mask_114,
  input        io_sc2mac_dat_mask_115,
  input        io_sc2mac_dat_mask_116,
  input        io_sc2mac_dat_mask_117,
  input        io_sc2mac_dat_mask_118,
  input        io_sc2mac_dat_mask_119,
  input        io_sc2mac_dat_mask_120,
  input        io_sc2mac_dat_mask_121,
  input        io_sc2mac_dat_mask_122,
  input        io_sc2mac_dat_mask_123,
  input        io_sc2mac_dat_mask_124,
  input        io_sc2mac_dat_mask_125,
  input        io_sc2mac_dat_mask_126,
  input        io_sc2mac_dat_mask_127,
  input  [8:0] io_sc2mac_dat_pd,
  input        io_sc2mac_dat_pvld,
  input  [7:0] io_sc2mac_wt_data_0,
  input  [7:0] io_sc2mac_wt_data_1,
  input  [7:0] io_sc2mac_wt_data_2,
  input  [7:0] io_sc2mac_wt_data_3,
  input  [7:0] io_sc2mac_wt_data_4,
  input  [7:0] io_sc2mac_wt_data_5,
  input  [7:0] io_sc2mac_wt_data_6,
  input  [7:0] io_sc2mac_wt_data_7,
  input  [7:0] io_sc2mac_wt_data_8,
  input  [7:0] io_sc2mac_wt_data_9,
  input  [7:0] io_sc2mac_wt_data_10,
  input  [7:0] io_sc2mac_wt_data_11,
  input  [7:0] io_sc2mac_wt_data_12,
  input  [7:0] io_sc2mac_wt_data_13,
  input  [7:0] io_sc2mac_wt_data_14,
  input  [7:0] io_sc2mac_wt_data_15,
  input  [7:0] io_sc2mac_wt_data_16,
  input  [7:0] io_sc2mac_wt_data_17,
  input  [7:0] io_sc2mac_wt_data_18,
  input  [7:0] io_sc2mac_wt_data_19,
  input  [7:0] io_sc2mac_wt_data_20,
  input  [7:0] io_sc2mac_wt_data_21,
  input  [7:0] io_sc2mac_wt_data_22,
  input  [7:0] io_sc2mac_wt_data_23,
  input  [7:0] io_sc2mac_wt_data_24,
  input  [7:0] io_sc2mac_wt_data_25,
  input  [7:0] io_sc2mac_wt_data_26,
  input  [7:0] io_sc2mac_wt_data_27,
  input  [7:0] io_sc2mac_wt_data_28,
  input  [7:0] io_sc2mac_wt_data_29,
  input  [7:0] io_sc2mac_wt_data_30,
  input  [7:0] io_sc2mac_wt_data_31,
  input  [7:0] io_sc2mac_wt_data_32,
  input  [7:0] io_sc2mac_wt_data_33,
  input  [7:0] io_sc2mac_wt_data_34,
  input  [7:0] io_sc2mac_wt_data_35,
  input  [7:0] io_sc2mac_wt_data_36,
  input  [7:0] io_sc2mac_wt_data_37,
  input  [7:0] io_sc2mac_wt_data_38,
  input  [7:0] io_sc2mac_wt_data_39,
  input  [7:0] io_sc2mac_wt_data_40,
  input  [7:0] io_sc2mac_wt_data_41,
  input  [7:0] io_sc2mac_wt_data_42,
  input  [7:0] io_sc2mac_wt_data_43,
  input  [7:0] io_sc2mac_wt_data_44,
  input  [7:0] io_sc2mac_wt_data_45,
  input  [7:0] io_sc2mac_wt_data_46,
  input  [7:0] io_sc2mac_wt_data_47,
  input  [7:0] io_sc2mac_wt_data_48,
  input  [7:0] io_sc2mac_wt_data_49,
  input  [7:0] io_sc2mac_wt_data_50,
  input  [7:0] io_sc2mac_wt_data_51,
  input  [7:0] io_sc2mac_wt_data_52,
  input  [7:0] io_sc2mac_wt_data_53,
  input  [7:0] io_sc2mac_wt_data_54,
  input  [7:0] io_sc2mac_wt_data_55,
  input  [7:0] io_sc2mac_wt_data_56,
  input  [7:0] io_sc2mac_wt_data_57,
  input  [7:0] io_sc2mac_wt_data_58,
  input  [7:0] io_sc2mac_wt_data_59,
  input  [7:0] io_sc2mac_wt_data_60,
  input  [7:0] io_sc2mac_wt_data_61,
  input  [7:0] io_sc2mac_wt_data_62,
  input  [7:0] io_sc2mac_wt_data_63,
  input  [7:0] io_sc2mac_wt_data_64,
  input  [7:0] io_sc2mac_wt_data_65,
  input  [7:0] io_sc2mac_wt_data_66,
  input  [7:0] io_sc2mac_wt_data_67,
  input  [7:0] io_sc2mac_wt_data_68,
  input  [7:0] io_sc2mac_wt_data_69,
  input  [7:0] io_sc2mac_wt_data_70,
  input  [7:0] io_sc2mac_wt_data_71,
  input  [7:0] io_sc2mac_wt_data_72,
  input  [7:0] io_sc2mac_wt_data_73,
  input  [7:0] io_sc2mac_wt_data_74,
  input  [7:0] io_sc2mac_wt_data_75,
  input  [7:0] io_sc2mac_wt_data_76,
  input  [7:0] io_sc2mac_wt_data_77,
  input  [7:0] io_sc2mac_wt_data_78,
  input  [7:0] io_sc2mac_wt_data_79,
  input  [7:0] io_sc2mac_wt_data_80,
  input  [7:0] io_sc2mac_wt_data_81,
  input  [7:0] io_sc2mac_wt_data_82,
  input  [7:0] io_sc2mac_wt_data_83,
  input  [7:0] io_sc2mac_wt_data_84,
  input  [7:0] io_sc2mac_wt_data_85,
  input  [7:0] io_sc2mac_wt_data_86,
  input  [7:0] io_sc2mac_wt_data_87,
  input  [7:0] io_sc2mac_wt_data_88,
  input  [7:0] io_sc2mac_wt_data_89,
  input  [7:0] io_sc2mac_wt_data_90,
  input  [7:0] io_sc2mac_wt_data_91,
  input  [7:0] io_sc2mac_wt_data_92,
  input  [7:0] io_sc2mac_wt_data_93,
  input  [7:0] io_sc2mac_wt_data_94,
  input  [7:0] io_sc2mac_wt_data_95,
  input  [7:0] io_sc2mac_wt_data_96,
  input  [7:0] io_sc2mac_wt_data_97,
  input  [7:0] io_sc2mac_wt_data_98,
  input  [7:0] io_sc2mac_wt_data_99,
  input  [7:0] io_sc2mac_wt_data_100,
  input  [7:0] io_sc2mac_wt_data_101,
  input  [7:0] io_sc2mac_wt_data_102,
  input  [7:0] io_sc2mac_wt_data_103,
  input  [7:0] io_sc2mac_wt_data_104,
  input  [7:0] io_sc2mac_wt_data_105,
  input  [7:0] io_sc2mac_wt_data_106,
  input  [7:0] io_sc2mac_wt_data_107,
  input  [7:0] io_sc2mac_wt_data_108,
  input  [7:0] io_sc2mac_wt_data_109,
  input  [7:0] io_sc2mac_wt_data_110,
  input  [7:0] io_sc2mac_wt_data_111,
  input  [7:0] io_sc2mac_wt_data_112,
  input  [7:0] io_sc2mac_wt_data_113,
  input  [7:0] io_sc2mac_wt_data_114,
  input  [7:0] io_sc2mac_wt_data_115,
  input  [7:0] io_sc2mac_wt_data_116,
  input  [7:0] io_sc2mac_wt_data_117,
  input  [7:0] io_sc2mac_wt_data_118,
  input  [7:0] io_sc2mac_wt_data_119,
  input  [7:0] io_sc2mac_wt_data_120,
  input  [7:0] io_sc2mac_wt_data_121,
  input  [7:0] io_sc2mac_wt_data_122,
  input  [7:0] io_sc2mac_wt_data_123,
  input  [7:0] io_sc2mac_wt_data_124,
  input  [7:0] io_sc2mac_wt_data_125,
  input  [7:0] io_sc2mac_wt_data_126,
  input  [7:0] io_sc2mac_wt_data_127,
  input        io_sc2mac_wt_mask_0,
  input        io_sc2mac_wt_mask_1,
  input        io_sc2mac_wt_mask_2,
  input        io_sc2mac_wt_mask_3,
  input        io_sc2mac_wt_mask_4,
  input        io_sc2mac_wt_mask_5,
  input        io_sc2mac_wt_mask_6,
  input        io_sc2mac_wt_mask_7,
  input        io_sc2mac_wt_mask_8,
  input        io_sc2mac_wt_mask_9,
  input        io_sc2mac_wt_mask_10,
  input        io_sc2mac_wt_mask_11,
  input        io_sc2mac_wt_mask_12,
  input        io_sc2mac_wt_mask_13,
  input        io_sc2mac_wt_mask_14,
  input        io_sc2mac_wt_mask_15,
  input        io_sc2mac_wt_mask_16,
  input        io_sc2mac_wt_mask_17,
  input        io_sc2mac_wt_mask_18,
  input        io_sc2mac_wt_mask_19,
  input        io_sc2mac_wt_mask_20,
  input        io_sc2mac_wt_mask_21,
  input        io_sc2mac_wt_mask_22,
  input        io_sc2mac_wt_mask_23,
  input        io_sc2mac_wt_mask_24,
  input        io_sc2mac_wt_mask_25,
  input        io_sc2mac_wt_mask_26,
  input        io_sc2mac_wt_mask_27,
  input        io_sc2mac_wt_mask_28,
  input        io_sc2mac_wt_mask_29,
  input        io_sc2mac_wt_mask_30,
  input        io_sc2mac_wt_mask_31,
  input        io_sc2mac_wt_mask_32,
  input        io_sc2mac_wt_mask_33,
  input        io_sc2mac_wt_mask_34,
  input        io_sc2mac_wt_mask_35,
  input        io_sc2mac_wt_mask_36,
  input        io_sc2mac_wt_mask_37,
  input        io_sc2mac_wt_mask_38,
  input        io_sc2mac_wt_mask_39,
  input        io_sc2mac_wt_mask_40,
  input        io_sc2mac_wt_mask_41,
  input        io_sc2mac_wt_mask_42,
  input        io_sc2mac_wt_mask_43,
  input        io_sc2mac_wt_mask_44,
  input        io_sc2mac_wt_mask_45,
  input        io_sc2mac_wt_mask_46,
  input        io_sc2mac_wt_mask_47,
  input        io_sc2mac_wt_mask_48,
  input        io_sc2mac_wt_mask_49,
  input        io_sc2mac_wt_mask_50,
  input        io_sc2mac_wt_mask_51,
  input        io_sc2mac_wt_mask_52,
  input        io_sc2mac_wt_mask_53,
  input        io_sc2mac_wt_mask_54,
  input        io_sc2mac_wt_mask_55,
  input        io_sc2mac_wt_mask_56,
  input        io_sc2mac_wt_mask_57,
  input        io_sc2mac_wt_mask_58,
  input        io_sc2mac_wt_mask_59,
  input        io_sc2mac_wt_mask_60,
  input        io_sc2mac_wt_mask_61,
  input        io_sc2mac_wt_mask_62,
  input        io_sc2mac_wt_mask_63,
  input        io_sc2mac_wt_mask_64,
  input        io_sc2mac_wt_mask_65,
  input        io_sc2mac_wt_mask_66,
  input        io_sc2mac_wt_mask_67,
  input        io_sc2mac_wt_mask_68,
  input        io_sc2mac_wt_mask_69,
  input        io_sc2mac_wt_mask_70,
  input        io_sc2mac_wt_mask_71,
  input        io_sc2mac_wt_mask_72,
  input        io_sc2mac_wt_mask_73,
  input        io_sc2mac_wt_mask_74,
  input        io_sc2mac_wt_mask_75,
  input        io_sc2mac_wt_mask_76,
  input        io_sc2mac_wt_mask_77,
  input        io_sc2mac_wt_mask_78,
  input        io_sc2mac_wt_mask_79,
  input        io_sc2mac_wt_mask_80,
  input        io_sc2mac_wt_mask_81,
  input        io_sc2mac_wt_mask_82,
  input        io_sc2mac_wt_mask_83,
  input        io_sc2mac_wt_mask_84,
  input        io_sc2mac_wt_mask_85,
  input        io_sc2mac_wt_mask_86,
  input        io_sc2mac_wt_mask_87,
  input        io_sc2mac_wt_mask_88,
  input        io_sc2mac_wt_mask_89,
  input        io_sc2mac_wt_mask_90,
  input        io_sc2mac_wt_mask_91,
  input        io_sc2mac_wt_mask_92,
  input        io_sc2mac_wt_mask_93,
  input        io_sc2mac_wt_mask_94,
  input        io_sc2mac_wt_mask_95,
  input        io_sc2mac_wt_mask_96,
  input        io_sc2mac_wt_mask_97,
  input        io_sc2mac_wt_mask_98,
  input        io_sc2mac_wt_mask_99,
  input        io_sc2mac_wt_mask_100,
  input        io_sc2mac_wt_mask_101,
  input        io_sc2mac_wt_mask_102,
  input        io_sc2mac_wt_mask_103,
  input        io_sc2mac_wt_mask_104,
  input        io_sc2mac_wt_mask_105,
  input        io_sc2mac_wt_mask_106,
  input        io_sc2mac_wt_mask_107,
  input        io_sc2mac_wt_mask_108,
  input        io_sc2mac_wt_mask_109,
  input        io_sc2mac_wt_mask_110,
  input        io_sc2mac_wt_mask_111,
  input        io_sc2mac_wt_mask_112,
  input        io_sc2mac_wt_mask_113,
  input        io_sc2mac_wt_mask_114,
  input        io_sc2mac_wt_mask_115,
  input        io_sc2mac_wt_mask_116,
  input        io_sc2mac_wt_mask_117,
  input        io_sc2mac_wt_mask_118,
  input        io_sc2mac_wt_mask_119,
  input        io_sc2mac_wt_mask_120,
  input        io_sc2mac_wt_mask_121,
  input        io_sc2mac_wt_mask_122,
  input        io_sc2mac_wt_mask_123,
  input        io_sc2mac_wt_mask_124,
  input        io_sc2mac_wt_mask_125,
  input        io_sc2mac_wt_mask_126,
  input        io_sc2mac_wt_mask_127,
  input        io_sc2mac_wt_sel_0,
  input        io_sc2mac_wt_pvld,
  output [7:0] io_in_dat_data_0,
  output [7:0] io_in_dat_data_1,
  output [7:0] io_in_dat_data_2,
  output [7:0] io_in_dat_data_3,
  output [7:0] io_in_dat_data_4,
  output [7:0] io_in_dat_data_5,
  output [7:0] io_in_dat_data_6,
  output [7:0] io_in_dat_data_7,
  output [7:0] io_in_dat_data_8,
  output [7:0] io_in_dat_data_9,
  output [7:0] io_in_dat_data_10,
  output [7:0] io_in_dat_data_11,
  output [7:0] io_in_dat_data_12,
  output [7:0] io_in_dat_data_13,
  output [7:0] io_in_dat_data_14,
  output [7:0] io_in_dat_data_15,
  output [7:0] io_in_dat_data_16,
  output [7:0] io_in_dat_data_17,
  output [7:0] io_in_dat_data_18,
  output [7:0] io_in_dat_data_19,
  output [7:0] io_in_dat_data_20,
  output [7:0] io_in_dat_data_21,
  output [7:0] io_in_dat_data_22,
  output [7:0] io_in_dat_data_23,
  output [7:0] io_in_dat_data_24,
  output [7:0] io_in_dat_data_25,
  output [7:0] io_in_dat_data_26,
  output [7:0] io_in_dat_data_27,
  output [7:0] io_in_dat_data_28,
  output [7:0] io_in_dat_data_29,
  output [7:0] io_in_dat_data_30,
  output [7:0] io_in_dat_data_31,
  output [7:0] io_in_dat_data_32,
  output [7:0] io_in_dat_data_33,
  output [7:0] io_in_dat_data_34,
  output [7:0] io_in_dat_data_35,
  output [7:0] io_in_dat_data_36,
  output [7:0] io_in_dat_data_37,
  output [7:0] io_in_dat_data_38,
  output [7:0] io_in_dat_data_39,
  output [7:0] io_in_dat_data_40,
  output [7:0] io_in_dat_data_41,
  output [7:0] io_in_dat_data_42,
  output [7:0] io_in_dat_data_43,
  output [7:0] io_in_dat_data_44,
  output [7:0] io_in_dat_data_45,
  output [7:0] io_in_dat_data_46,
  output [7:0] io_in_dat_data_47,
  output [7:0] io_in_dat_data_48,
  output [7:0] io_in_dat_data_49,
  output [7:0] io_in_dat_data_50,
  output [7:0] io_in_dat_data_51,
  output [7:0] io_in_dat_data_52,
  output [7:0] io_in_dat_data_53,
  output [7:0] io_in_dat_data_54,
  output [7:0] io_in_dat_data_55,
  output [7:0] io_in_dat_data_56,
  output [7:0] io_in_dat_data_57,
  output [7:0] io_in_dat_data_58,
  output [7:0] io_in_dat_data_59,
  output [7:0] io_in_dat_data_60,
  output [7:0] io_in_dat_data_61,
  output [7:0] io_in_dat_data_62,
  output [7:0] io_in_dat_data_63,
  output [7:0] io_in_dat_data_64,
  output [7:0] io_in_dat_data_65,
  output [7:0] io_in_dat_data_66,
  output [7:0] io_in_dat_data_67,
  output [7:0] io_in_dat_data_68,
  output [7:0] io_in_dat_data_69,
  output [7:0] io_in_dat_data_70,
  output [7:0] io_in_dat_data_71,
  output [7:0] io_in_dat_data_72,
  output [7:0] io_in_dat_data_73,
  output [7:0] io_in_dat_data_74,
  output [7:0] io_in_dat_data_75,
  output [7:0] io_in_dat_data_76,
  output [7:0] io_in_dat_data_77,
  output [7:0] io_in_dat_data_78,
  output [7:0] io_in_dat_data_79,
  output [7:0] io_in_dat_data_80,
  output [7:0] io_in_dat_data_81,
  output [7:0] io_in_dat_data_82,
  output [7:0] io_in_dat_data_83,
  output [7:0] io_in_dat_data_84,
  output [7:0] io_in_dat_data_85,
  output [7:0] io_in_dat_data_86,
  output [7:0] io_in_dat_data_87,
  output [7:0] io_in_dat_data_88,
  output [7:0] io_in_dat_data_89,
  output [7:0] io_in_dat_data_90,
  output [7:0] io_in_dat_data_91,
  output [7:0] io_in_dat_data_92,
  output [7:0] io_in_dat_data_93,
  output [7:0] io_in_dat_data_94,
  output [7:0] io_in_dat_data_95,
  output [7:0] io_in_dat_data_96,
  output [7:0] io_in_dat_data_97,
  output [7:0] io_in_dat_data_98,
  output [7:0] io_in_dat_data_99,
  output [7:0] io_in_dat_data_100,
  output [7:0] io_in_dat_data_101,
  output [7:0] io_in_dat_data_102,
  output [7:0] io_in_dat_data_103,
  output [7:0] io_in_dat_data_104,
  output [7:0] io_in_dat_data_105,
  output [7:0] io_in_dat_data_106,
  output [7:0] io_in_dat_data_107,
  output [7:0] io_in_dat_data_108,
  output [7:0] io_in_dat_data_109,
  output [7:0] io_in_dat_data_110,
  output [7:0] io_in_dat_data_111,
  output [7:0] io_in_dat_data_112,
  output [7:0] io_in_dat_data_113,
  output [7:0] io_in_dat_data_114,
  output [7:0] io_in_dat_data_115,
  output [7:0] io_in_dat_data_116,
  output [7:0] io_in_dat_data_117,
  output [7:0] io_in_dat_data_118,
  output [7:0] io_in_dat_data_119,
  output [7:0] io_in_dat_data_120,
  output [7:0] io_in_dat_data_121,
  output [7:0] io_in_dat_data_122,
  output [7:0] io_in_dat_data_123,
  output [7:0] io_in_dat_data_124,
  output [7:0] io_in_dat_data_125,
  output [7:0] io_in_dat_data_126,
  output [7:0] io_in_dat_data_127,
  output       io_in_dat_mask_0,
  output       io_in_dat_mask_1,
  output       io_in_dat_mask_2,
  output       io_in_dat_mask_3,
  output       io_in_dat_mask_4,
  output       io_in_dat_mask_5,
  output       io_in_dat_mask_6,
  output       io_in_dat_mask_7,
  output       io_in_dat_mask_8,
  output       io_in_dat_mask_9,
  output       io_in_dat_mask_10,
  output       io_in_dat_mask_11,
  output       io_in_dat_mask_12,
  output       io_in_dat_mask_13,
  output       io_in_dat_mask_14,
  output       io_in_dat_mask_15,
  output       io_in_dat_mask_16,
  output       io_in_dat_mask_17,
  output       io_in_dat_mask_18,
  output       io_in_dat_mask_19,
  output       io_in_dat_mask_20,
  output       io_in_dat_mask_21,
  output       io_in_dat_mask_22,
  output       io_in_dat_mask_23,
  output       io_in_dat_mask_24,
  output       io_in_dat_mask_25,
  output       io_in_dat_mask_26,
  output       io_in_dat_mask_27,
  output       io_in_dat_mask_28,
  output       io_in_dat_mask_29,
  output       io_in_dat_mask_30,
  output       io_in_dat_mask_31,
  output       io_in_dat_mask_32,
  output       io_in_dat_mask_33,
  output       io_in_dat_mask_34,
  output       io_in_dat_mask_35,
  output       io_in_dat_mask_36,
  output       io_in_dat_mask_37,
  output       io_in_dat_mask_38,
  output       io_in_dat_mask_39,
  output       io_in_dat_mask_40,
  output       io_in_dat_mask_41,
  output       io_in_dat_mask_42,
  output       io_in_dat_mask_43,
  output       io_in_dat_mask_44,
  output       io_in_dat_mask_45,
  output       io_in_dat_mask_46,
  output       io_in_dat_mask_47,
  output       io_in_dat_mask_48,
  output       io_in_dat_mask_49,
  output       io_in_dat_mask_50,
  output       io_in_dat_mask_51,
  output       io_in_dat_mask_52,
  output       io_in_dat_mask_53,
  output       io_in_dat_mask_54,
  output       io_in_dat_mask_55,
  output       io_in_dat_mask_56,
  output       io_in_dat_mask_57,
  output       io_in_dat_mask_58,
  output       io_in_dat_mask_59,
  output       io_in_dat_mask_60,
  output       io_in_dat_mask_61,
  output       io_in_dat_mask_62,
  output       io_in_dat_mask_63,
  output       io_in_dat_mask_64,
  output       io_in_dat_mask_65,
  output       io_in_dat_mask_66,
  output       io_in_dat_mask_67,
  output       io_in_dat_mask_68,
  output       io_in_dat_mask_69,
  output       io_in_dat_mask_70,
  output       io_in_dat_mask_71,
  output       io_in_dat_mask_72,
  output       io_in_dat_mask_73,
  output       io_in_dat_mask_74,
  output       io_in_dat_mask_75,
  output       io_in_dat_mask_76,
  output       io_in_dat_mask_77,
  output       io_in_dat_mask_78,
  output       io_in_dat_mask_79,
  output       io_in_dat_mask_80,
  output       io_in_dat_mask_81,
  output       io_in_dat_mask_82,
  output       io_in_dat_mask_83,
  output       io_in_dat_mask_84,
  output       io_in_dat_mask_85,
  output       io_in_dat_mask_86,
  output       io_in_dat_mask_87,
  output       io_in_dat_mask_88,
  output       io_in_dat_mask_89,
  output       io_in_dat_mask_90,
  output       io_in_dat_mask_91,
  output       io_in_dat_mask_92,
  output       io_in_dat_mask_93,
  output       io_in_dat_mask_94,
  output       io_in_dat_mask_95,
  output       io_in_dat_mask_96,
  output       io_in_dat_mask_97,
  output       io_in_dat_mask_98,
  output       io_in_dat_mask_99,
  output       io_in_dat_mask_100,
  output       io_in_dat_mask_101,
  output       io_in_dat_mask_102,
  output       io_in_dat_mask_103,
  output       io_in_dat_mask_104,
  output       io_in_dat_mask_105,
  output       io_in_dat_mask_106,
  output       io_in_dat_mask_107,
  output       io_in_dat_mask_108,
  output       io_in_dat_mask_109,
  output       io_in_dat_mask_110,
  output       io_in_dat_mask_111,
  output       io_in_dat_mask_112,
  output       io_in_dat_mask_113,
  output       io_in_dat_mask_114,
  output       io_in_dat_mask_115,
  output       io_in_dat_mask_116,
  output       io_in_dat_mask_117,
  output       io_in_dat_mask_118,
  output       io_in_dat_mask_119,
  output       io_in_dat_mask_120,
  output       io_in_dat_mask_121,
  output       io_in_dat_mask_122,
  output       io_in_dat_mask_123,
  output       io_in_dat_mask_124,
  output       io_in_dat_mask_125,
  output       io_in_dat_mask_126,
  output       io_in_dat_mask_127,
  output [8:0] io_in_dat_pd,
  output       io_in_dat_pvld,
  output       io_in_dat_stripe_st,
  output       io_in_dat_stripe_end,
  output [7:0] io_in_wt_data_0,
  output [7:0] io_in_wt_data_1,
  output [7:0] io_in_wt_data_2,
  output [7:0] io_in_wt_data_3,
  output [7:0] io_in_wt_data_4,
  output [7:0] io_in_wt_data_5,
  output [7:0] io_in_wt_data_6,
  output [7:0] io_in_wt_data_7,
  output [7:0] io_in_wt_data_8,
  output [7:0] io_in_wt_data_9,
  output [7:0] io_in_wt_data_10,
  output [7:0] io_in_wt_data_11,
  output [7:0] io_in_wt_data_12,
  output [7:0] io_in_wt_data_13,
  output [7:0] io_in_wt_data_14,
  output [7:0] io_in_wt_data_15,
  output [7:0] io_in_wt_data_16,
  output [7:0] io_in_wt_data_17,
  output [7:0] io_in_wt_data_18,
  output [7:0] io_in_wt_data_19,
  output [7:0] io_in_wt_data_20,
  output [7:0] io_in_wt_data_21,
  output [7:0] io_in_wt_data_22,
  output [7:0] io_in_wt_data_23,
  output [7:0] io_in_wt_data_24,
  output [7:0] io_in_wt_data_25,
  output [7:0] io_in_wt_data_26,
  output [7:0] io_in_wt_data_27,
  output [7:0] io_in_wt_data_28,
  output [7:0] io_in_wt_data_29,
  output [7:0] io_in_wt_data_30,
  output [7:0] io_in_wt_data_31,
  output [7:0] io_in_wt_data_32,
  output [7:0] io_in_wt_data_33,
  output [7:0] io_in_wt_data_34,
  output [7:0] io_in_wt_data_35,
  output [7:0] io_in_wt_data_36,
  output [7:0] io_in_wt_data_37,
  output [7:0] io_in_wt_data_38,
  output [7:0] io_in_wt_data_39,
  output [7:0] io_in_wt_data_40,
  output [7:0] io_in_wt_data_41,
  output [7:0] io_in_wt_data_42,
  output [7:0] io_in_wt_data_43,
  output [7:0] io_in_wt_data_44,
  output [7:0] io_in_wt_data_45,
  output [7:0] io_in_wt_data_46,
  output [7:0] io_in_wt_data_47,
  output [7:0] io_in_wt_data_48,
  output [7:0] io_in_wt_data_49,
  output [7:0] io_in_wt_data_50,
  output [7:0] io_in_wt_data_51,
  output [7:0] io_in_wt_data_52,
  output [7:0] io_in_wt_data_53,
  output [7:0] io_in_wt_data_54,
  output [7:0] io_in_wt_data_55,
  output [7:0] io_in_wt_data_56,
  output [7:0] io_in_wt_data_57,
  output [7:0] io_in_wt_data_58,
  output [7:0] io_in_wt_data_59,
  output [7:0] io_in_wt_data_60,
  output [7:0] io_in_wt_data_61,
  output [7:0] io_in_wt_data_62,
  output [7:0] io_in_wt_data_63,
  output [7:0] io_in_wt_data_64,
  output [7:0] io_in_wt_data_65,
  output [7:0] io_in_wt_data_66,
  output [7:0] io_in_wt_data_67,
  output [7:0] io_in_wt_data_68,
  output [7:0] io_in_wt_data_69,
  output [7:0] io_in_wt_data_70,
  output [7:0] io_in_wt_data_71,
  output [7:0] io_in_wt_data_72,
  output [7:0] io_in_wt_data_73,
  output [7:0] io_in_wt_data_74,
  output [7:0] io_in_wt_data_75,
  output [7:0] io_in_wt_data_76,
  output [7:0] io_in_wt_data_77,
  output [7:0] io_in_wt_data_78,
  output [7:0] io_in_wt_data_79,
  output [7:0] io_in_wt_data_80,
  output [7:0] io_in_wt_data_81,
  output [7:0] io_in_wt_data_82,
  output [7:0] io_in_wt_data_83,
  output [7:0] io_in_wt_data_84,
  output [7:0] io_in_wt_data_85,
  output [7:0] io_in_wt_data_86,
  output [7:0] io_in_wt_data_87,
  output [7:0] io_in_wt_data_88,
  output [7:0] io_in_wt_data_89,
  output [7:0] io_in_wt_data_90,
  output [7:0] io_in_wt_data_91,
  output [7:0] io_in_wt_data_92,
  output [7:0] io_in_wt_data_93,
  output [7:0] io_in_wt_data_94,
  output [7:0] io_in_wt_data_95,
  output [7:0] io_in_wt_data_96,
  output [7:0] io_in_wt_data_97,
  output [7:0] io_in_wt_data_98,
  output [7:0] io_in_wt_data_99,
  output [7:0] io_in_wt_data_100,
  output [7:0] io_in_wt_data_101,
  output [7:0] io_in_wt_data_102,
  output [7:0] io_in_wt_data_103,
  output [7:0] io_in_wt_data_104,
  output [7:0] io_in_wt_data_105,
  output [7:0] io_in_wt_data_106,
  output [7:0] io_in_wt_data_107,
  output [7:0] io_in_wt_data_108,
  output [7:0] io_in_wt_data_109,
  output [7:0] io_in_wt_data_110,
  output [7:0] io_in_wt_data_111,
  output [7:0] io_in_wt_data_112,
  output [7:0] io_in_wt_data_113,
  output [7:0] io_in_wt_data_114,
  output [7:0] io_in_wt_data_115,
  output [7:0] io_in_wt_data_116,
  output [7:0] io_in_wt_data_117,
  output [7:0] io_in_wt_data_118,
  output [7:0] io_in_wt_data_119,
  output [7:0] io_in_wt_data_120,
  output [7:0] io_in_wt_data_121,
  output [7:0] io_in_wt_data_122,
  output [7:0] io_in_wt_data_123,
  output [7:0] io_in_wt_data_124,
  output [7:0] io_in_wt_data_125,
  output [7:0] io_in_wt_data_126,
  output [7:0] io_in_wt_data_127,
  output       io_in_wt_mask_0,
  output       io_in_wt_mask_1,
  output       io_in_wt_mask_2,
  output       io_in_wt_mask_3,
  output       io_in_wt_mask_4,
  output       io_in_wt_mask_5,
  output       io_in_wt_mask_6,
  output       io_in_wt_mask_7,
  output       io_in_wt_mask_8,
  output       io_in_wt_mask_9,
  output       io_in_wt_mask_10,
  output       io_in_wt_mask_11,
  output       io_in_wt_mask_12,
  output       io_in_wt_mask_13,
  output       io_in_wt_mask_14,
  output       io_in_wt_mask_15,
  output       io_in_wt_mask_16,
  output       io_in_wt_mask_17,
  output       io_in_wt_mask_18,
  output       io_in_wt_mask_19,
  output       io_in_wt_mask_20,
  output       io_in_wt_mask_21,
  output       io_in_wt_mask_22,
  output       io_in_wt_mask_23,
  output       io_in_wt_mask_24,
  output       io_in_wt_mask_25,
  output       io_in_wt_mask_26,
  output       io_in_wt_mask_27,
  output       io_in_wt_mask_28,
  output       io_in_wt_mask_29,
  output       io_in_wt_mask_30,
  output       io_in_wt_mask_31,
  output       io_in_wt_mask_32,
  output       io_in_wt_mask_33,
  output       io_in_wt_mask_34,
  output       io_in_wt_mask_35,
  output       io_in_wt_mask_36,
  output       io_in_wt_mask_37,
  output       io_in_wt_mask_38,
  output       io_in_wt_mask_39,
  output       io_in_wt_mask_40,
  output       io_in_wt_mask_41,
  output       io_in_wt_mask_42,
  output       io_in_wt_mask_43,
  output       io_in_wt_mask_44,
  output       io_in_wt_mask_45,
  output       io_in_wt_mask_46,
  output       io_in_wt_mask_47,
  output       io_in_wt_mask_48,
  output       io_in_wt_mask_49,
  output       io_in_wt_mask_50,
  output       io_in_wt_mask_51,
  output       io_in_wt_mask_52,
  output       io_in_wt_mask_53,
  output       io_in_wt_mask_54,
  output       io_in_wt_mask_55,
  output       io_in_wt_mask_56,
  output       io_in_wt_mask_57,
  output       io_in_wt_mask_58,
  output       io_in_wt_mask_59,
  output       io_in_wt_mask_60,
  output       io_in_wt_mask_61,
  output       io_in_wt_mask_62,
  output       io_in_wt_mask_63,
  output       io_in_wt_mask_64,
  output       io_in_wt_mask_65,
  output       io_in_wt_mask_66,
  output       io_in_wt_mask_67,
  output       io_in_wt_mask_68,
  output       io_in_wt_mask_69,
  output       io_in_wt_mask_70,
  output       io_in_wt_mask_71,
  output       io_in_wt_mask_72,
  output       io_in_wt_mask_73,
  output       io_in_wt_mask_74,
  output       io_in_wt_mask_75,
  output       io_in_wt_mask_76,
  output       io_in_wt_mask_77,
  output       io_in_wt_mask_78,
  output       io_in_wt_mask_79,
  output       io_in_wt_mask_80,
  output       io_in_wt_mask_81,
  output       io_in_wt_mask_82,
  output       io_in_wt_mask_83,
  output       io_in_wt_mask_84,
  output       io_in_wt_mask_85,
  output       io_in_wt_mask_86,
  output       io_in_wt_mask_87,
  output       io_in_wt_mask_88,
  output       io_in_wt_mask_89,
  output       io_in_wt_mask_90,
  output       io_in_wt_mask_91,
  output       io_in_wt_mask_92,
  output       io_in_wt_mask_93,
  output       io_in_wt_mask_94,
  output       io_in_wt_mask_95,
  output       io_in_wt_mask_96,
  output       io_in_wt_mask_97,
  output       io_in_wt_mask_98,
  output       io_in_wt_mask_99,
  output       io_in_wt_mask_100,
  output       io_in_wt_mask_101,
  output       io_in_wt_mask_102,
  output       io_in_wt_mask_103,
  output       io_in_wt_mask_104,
  output       io_in_wt_mask_105,
  output       io_in_wt_mask_106,
  output       io_in_wt_mask_107,
  output       io_in_wt_mask_108,
  output       io_in_wt_mask_109,
  output       io_in_wt_mask_110,
  output       io_in_wt_mask_111,
  output       io_in_wt_mask_112,
  output       io_in_wt_mask_113,
  output       io_in_wt_mask_114,
  output       io_in_wt_mask_115,
  output       io_in_wt_mask_116,
  output       io_in_wt_mask_117,
  output       io_in_wt_mask_118,
  output       io_in_wt_mask_119,
  output       io_in_wt_mask_120,
  output       io_in_wt_mask_121,
  output       io_in_wt_mask_122,
  output       io_in_wt_mask_123,
  output       io_in_wt_mask_124,
  output       io_in_wt_mask_125,
  output       io_in_wt_mask_126,
  output       io_in_wt_mask_127,
  output       io_in_wt_sel_0,
  output       io_in_wt_pvld
);
  reg [7:0] in_rt_dat_data_d_1_0; // @[retiming.scala 9:92]
  reg [31:0] _RAND_0;
  reg [7:0] in_rt_dat_data_d_1_1; // @[retiming.scala 9:92]
  reg [31:0] _RAND_1;
  reg [7:0] in_rt_dat_data_d_1_2; // @[retiming.scala 9:92]
  reg [31:0] _RAND_2;
  reg [7:0] in_rt_dat_data_d_1_3; // @[retiming.scala 9:92]
  reg [31:0] _RAND_3;
  reg [7:0] in_rt_dat_data_d_1_4; // @[retiming.scala 9:92]
  reg [31:0] _RAND_4;
  reg [7:0] in_rt_dat_data_d_1_5; // @[retiming.scala 9:92]
  reg [31:0] _RAND_5;
  reg [7:0] in_rt_dat_data_d_1_6; // @[retiming.scala 9:92]
  reg [31:0] _RAND_6;
  reg [7:0] in_rt_dat_data_d_1_7; // @[retiming.scala 9:92]
  reg [31:0] _RAND_7;
  reg [7:0] in_rt_dat_data_d_1_8; // @[retiming.scala 9:92]
  reg [31:0] _RAND_8;
  reg [7:0] in_rt_dat_data_d_1_9; // @[retiming.scala 9:92]
  reg [31:0] _RAND_9;
  reg [7:0] in_rt_dat_data_d_1_10; // @[retiming.scala 9:92]
  reg [31:0] _RAND_10;
  reg [7:0] in_rt_dat_data_d_1_11; // @[retiming.scala 9:92]
  reg [31:0] _RAND_11;
  reg [7:0] in_rt_dat_data_d_1_12; // @[retiming.scala 9:92]
  reg [31:0] _RAND_12;
  reg [7:0] in_rt_dat_data_d_1_13; // @[retiming.scala 9:92]
  reg [31:0] _RAND_13;
  reg [7:0] in_rt_dat_data_d_1_14; // @[retiming.scala 9:92]
  reg [31:0] _RAND_14;
  reg [7:0] in_rt_dat_data_d_1_15; // @[retiming.scala 9:92]
  reg [31:0] _RAND_15;
  reg [7:0] in_rt_dat_data_d_1_16; // @[retiming.scala 9:92]
  reg [31:0] _RAND_16;
  reg [7:0] in_rt_dat_data_d_1_17; // @[retiming.scala 9:92]
  reg [31:0] _RAND_17;
  reg [7:0] in_rt_dat_data_d_1_18; // @[retiming.scala 9:92]
  reg [31:0] _RAND_18;
  reg [7:0] in_rt_dat_data_d_1_19; // @[retiming.scala 9:92]
  reg [31:0] _RAND_19;
  reg [7:0] in_rt_dat_data_d_1_20; // @[retiming.scala 9:92]
  reg [31:0] _RAND_20;
  reg [7:0] in_rt_dat_data_d_1_21; // @[retiming.scala 9:92]
  reg [31:0] _RAND_21;
  reg [7:0] in_rt_dat_data_d_1_22; // @[retiming.scala 9:92]
  reg [31:0] _RAND_22;
  reg [7:0] in_rt_dat_data_d_1_23; // @[retiming.scala 9:92]
  reg [31:0] _RAND_23;
  reg [7:0] in_rt_dat_data_d_1_24; // @[retiming.scala 9:92]
  reg [31:0] _RAND_24;
  reg [7:0] in_rt_dat_data_d_1_25; // @[retiming.scala 9:92]
  reg [31:0] _RAND_25;
  reg [7:0] in_rt_dat_data_d_1_26; // @[retiming.scala 9:92]
  reg [31:0] _RAND_26;
  reg [7:0] in_rt_dat_data_d_1_27; // @[retiming.scala 9:92]
  reg [31:0] _RAND_27;
  reg [7:0] in_rt_dat_data_d_1_28; // @[retiming.scala 9:92]
  reg [31:0] _RAND_28;
  reg [7:0] in_rt_dat_data_d_1_29; // @[retiming.scala 9:92]
  reg [31:0] _RAND_29;
  reg [7:0] in_rt_dat_data_d_1_30; // @[retiming.scala 9:92]
  reg [31:0] _RAND_30;
  reg [7:0] in_rt_dat_data_d_1_31; // @[retiming.scala 9:92]
  reg [31:0] _RAND_31;
  reg [7:0] in_rt_dat_data_d_1_32; // @[retiming.scala 9:92]
  reg [31:0] _RAND_32;
  reg [7:0] in_rt_dat_data_d_1_33; // @[retiming.scala 9:92]
  reg [31:0] _RAND_33;
  reg [7:0] in_rt_dat_data_d_1_34; // @[retiming.scala 9:92]
  reg [31:0] _RAND_34;
  reg [7:0] in_rt_dat_data_d_1_35; // @[retiming.scala 9:92]
  reg [31:0] _RAND_35;
  reg [7:0] in_rt_dat_data_d_1_36; // @[retiming.scala 9:92]
  reg [31:0] _RAND_36;
  reg [7:0] in_rt_dat_data_d_1_37; // @[retiming.scala 9:92]
  reg [31:0] _RAND_37;
  reg [7:0] in_rt_dat_data_d_1_38; // @[retiming.scala 9:92]
  reg [31:0] _RAND_38;
  reg [7:0] in_rt_dat_data_d_1_39; // @[retiming.scala 9:92]
  reg [31:0] _RAND_39;
  reg [7:0] in_rt_dat_data_d_1_40; // @[retiming.scala 9:92]
  reg [31:0] _RAND_40;
  reg [7:0] in_rt_dat_data_d_1_41; // @[retiming.scala 9:92]
  reg [31:0] _RAND_41;
  reg [7:0] in_rt_dat_data_d_1_42; // @[retiming.scala 9:92]
  reg [31:0] _RAND_42;
  reg [7:0] in_rt_dat_data_d_1_43; // @[retiming.scala 9:92]
  reg [31:0] _RAND_43;
  reg [7:0] in_rt_dat_data_d_1_44; // @[retiming.scala 9:92]
  reg [31:0] _RAND_44;
  reg [7:0] in_rt_dat_data_d_1_45; // @[retiming.scala 9:92]
  reg [31:0] _RAND_45;
  reg [7:0] in_rt_dat_data_d_1_46; // @[retiming.scala 9:92]
  reg [31:0] _RAND_46;
  reg [7:0] in_rt_dat_data_d_1_47; // @[retiming.scala 9:92]
  reg [31:0] _RAND_47;
  reg [7:0] in_rt_dat_data_d_1_48; // @[retiming.scala 9:92]
  reg [31:0] _RAND_48;
  reg [7:0] in_rt_dat_data_d_1_49; // @[retiming.scala 9:92]
  reg [31:0] _RAND_49;
  reg [7:0] in_rt_dat_data_d_1_50; // @[retiming.scala 9:92]
  reg [31:0] _RAND_50;
  reg [7:0] in_rt_dat_data_d_1_51; // @[retiming.scala 9:92]
  reg [31:0] _RAND_51;
  reg [7:0] in_rt_dat_data_d_1_52; // @[retiming.scala 9:92]
  reg [31:0] _RAND_52;
  reg [7:0] in_rt_dat_data_d_1_53; // @[retiming.scala 9:92]
  reg [31:0] _RAND_53;
  reg [7:0] in_rt_dat_data_d_1_54; // @[retiming.scala 9:92]
  reg [31:0] _RAND_54;
  reg [7:0] in_rt_dat_data_d_1_55; // @[retiming.scala 9:92]
  reg [31:0] _RAND_55;
  reg [7:0] in_rt_dat_data_d_1_56; // @[retiming.scala 9:92]
  reg [31:0] _RAND_56;
  reg [7:0] in_rt_dat_data_d_1_57; // @[retiming.scala 9:92]
  reg [31:0] _RAND_57;
  reg [7:0] in_rt_dat_data_d_1_58; // @[retiming.scala 9:92]
  reg [31:0] _RAND_58;
  reg [7:0] in_rt_dat_data_d_1_59; // @[retiming.scala 9:92]
  reg [31:0] _RAND_59;
  reg [7:0] in_rt_dat_data_d_1_60; // @[retiming.scala 9:92]
  reg [31:0] _RAND_60;
  reg [7:0] in_rt_dat_data_d_1_61; // @[retiming.scala 9:92]
  reg [31:0] _RAND_61;
  reg [7:0] in_rt_dat_data_d_1_62; // @[retiming.scala 9:92]
  reg [31:0] _RAND_62;
  reg [7:0] in_rt_dat_data_d_1_63; // @[retiming.scala 9:92]
  reg [31:0] _RAND_63;
  reg [7:0] in_rt_dat_data_d_1_64; // @[retiming.scala 9:92]
  reg [31:0] _RAND_64;
  reg [7:0] in_rt_dat_data_d_1_65; // @[retiming.scala 9:92]
  reg [31:0] _RAND_65;
  reg [7:0] in_rt_dat_data_d_1_66; // @[retiming.scala 9:92]
  reg [31:0] _RAND_66;
  reg [7:0] in_rt_dat_data_d_1_67; // @[retiming.scala 9:92]
  reg [31:0] _RAND_67;
  reg [7:0] in_rt_dat_data_d_1_68; // @[retiming.scala 9:92]
  reg [31:0] _RAND_68;
  reg [7:0] in_rt_dat_data_d_1_69; // @[retiming.scala 9:92]
  reg [31:0] _RAND_69;
  reg [7:0] in_rt_dat_data_d_1_70; // @[retiming.scala 9:92]
  reg [31:0] _RAND_70;
  reg [7:0] in_rt_dat_data_d_1_71; // @[retiming.scala 9:92]
  reg [31:0] _RAND_71;
  reg [7:0] in_rt_dat_data_d_1_72; // @[retiming.scala 9:92]
  reg [31:0] _RAND_72;
  reg [7:0] in_rt_dat_data_d_1_73; // @[retiming.scala 9:92]
  reg [31:0] _RAND_73;
  reg [7:0] in_rt_dat_data_d_1_74; // @[retiming.scala 9:92]
  reg [31:0] _RAND_74;
  reg [7:0] in_rt_dat_data_d_1_75; // @[retiming.scala 9:92]
  reg [31:0] _RAND_75;
  reg [7:0] in_rt_dat_data_d_1_76; // @[retiming.scala 9:92]
  reg [31:0] _RAND_76;
  reg [7:0] in_rt_dat_data_d_1_77; // @[retiming.scala 9:92]
  reg [31:0] _RAND_77;
  reg [7:0] in_rt_dat_data_d_1_78; // @[retiming.scala 9:92]
  reg [31:0] _RAND_78;
  reg [7:0] in_rt_dat_data_d_1_79; // @[retiming.scala 9:92]
  reg [31:0] _RAND_79;
  reg [7:0] in_rt_dat_data_d_1_80; // @[retiming.scala 9:92]
  reg [31:0] _RAND_80;
  reg [7:0] in_rt_dat_data_d_1_81; // @[retiming.scala 9:92]
  reg [31:0] _RAND_81;
  reg [7:0] in_rt_dat_data_d_1_82; // @[retiming.scala 9:92]
  reg [31:0] _RAND_82;
  reg [7:0] in_rt_dat_data_d_1_83; // @[retiming.scala 9:92]
  reg [31:0] _RAND_83;
  reg [7:0] in_rt_dat_data_d_1_84; // @[retiming.scala 9:92]
  reg [31:0] _RAND_84;
  reg [7:0] in_rt_dat_data_d_1_85; // @[retiming.scala 9:92]
  reg [31:0] _RAND_85;
  reg [7:0] in_rt_dat_data_d_1_86; // @[retiming.scala 9:92]
  reg [31:0] _RAND_86;
  reg [7:0] in_rt_dat_data_d_1_87; // @[retiming.scala 9:92]
  reg [31:0] _RAND_87;
  reg [7:0] in_rt_dat_data_d_1_88; // @[retiming.scala 9:92]
  reg [31:0] _RAND_88;
  reg [7:0] in_rt_dat_data_d_1_89; // @[retiming.scala 9:92]
  reg [31:0] _RAND_89;
  reg [7:0] in_rt_dat_data_d_1_90; // @[retiming.scala 9:92]
  reg [31:0] _RAND_90;
  reg [7:0] in_rt_dat_data_d_1_91; // @[retiming.scala 9:92]
  reg [31:0] _RAND_91;
  reg [7:0] in_rt_dat_data_d_1_92; // @[retiming.scala 9:92]
  reg [31:0] _RAND_92;
  reg [7:0] in_rt_dat_data_d_1_93; // @[retiming.scala 9:92]
  reg [31:0] _RAND_93;
  reg [7:0] in_rt_dat_data_d_1_94; // @[retiming.scala 9:92]
  reg [31:0] _RAND_94;
  reg [7:0] in_rt_dat_data_d_1_95; // @[retiming.scala 9:92]
  reg [31:0] _RAND_95;
  reg [7:0] in_rt_dat_data_d_1_96; // @[retiming.scala 9:92]
  reg [31:0] _RAND_96;
  reg [7:0] in_rt_dat_data_d_1_97; // @[retiming.scala 9:92]
  reg [31:0] _RAND_97;
  reg [7:0] in_rt_dat_data_d_1_98; // @[retiming.scala 9:92]
  reg [31:0] _RAND_98;
  reg [7:0] in_rt_dat_data_d_1_99; // @[retiming.scala 9:92]
  reg [31:0] _RAND_99;
  reg [7:0] in_rt_dat_data_d_1_100; // @[retiming.scala 9:92]
  reg [31:0] _RAND_100;
  reg [7:0] in_rt_dat_data_d_1_101; // @[retiming.scala 9:92]
  reg [31:0] _RAND_101;
  reg [7:0] in_rt_dat_data_d_1_102; // @[retiming.scala 9:92]
  reg [31:0] _RAND_102;
  reg [7:0] in_rt_dat_data_d_1_103; // @[retiming.scala 9:92]
  reg [31:0] _RAND_103;
  reg [7:0] in_rt_dat_data_d_1_104; // @[retiming.scala 9:92]
  reg [31:0] _RAND_104;
  reg [7:0] in_rt_dat_data_d_1_105; // @[retiming.scala 9:92]
  reg [31:0] _RAND_105;
  reg [7:0] in_rt_dat_data_d_1_106; // @[retiming.scala 9:92]
  reg [31:0] _RAND_106;
  reg [7:0] in_rt_dat_data_d_1_107; // @[retiming.scala 9:92]
  reg [31:0] _RAND_107;
  reg [7:0] in_rt_dat_data_d_1_108; // @[retiming.scala 9:92]
  reg [31:0] _RAND_108;
  reg [7:0] in_rt_dat_data_d_1_109; // @[retiming.scala 9:92]
  reg [31:0] _RAND_109;
  reg [7:0] in_rt_dat_data_d_1_110; // @[retiming.scala 9:92]
  reg [31:0] _RAND_110;
  reg [7:0] in_rt_dat_data_d_1_111; // @[retiming.scala 9:92]
  reg [31:0] _RAND_111;
  reg [7:0] in_rt_dat_data_d_1_112; // @[retiming.scala 9:92]
  reg [31:0] _RAND_112;
  reg [7:0] in_rt_dat_data_d_1_113; // @[retiming.scala 9:92]
  reg [31:0] _RAND_113;
  reg [7:0] in_rt_dat_data_d_1_114; // @[retiming.scala 9:92]
  reg [31:0] _RAND_114;
  reg [7:0] in_rt_dat_data_d_1_115; // @[retiming.scala 9:92]
  reg [31:0] _RAND_115;
  reg [7:0] in_rt_dat_data_d_1_116; // @[retiming.scala 9:92]
  reg [31:0] _RAND_116;
  reg [7:0] in_rt_dat_data_d_1_117; // @[retiming.scala 9:92]
  reg [31:0] _RAND_117;
  reg [7:0] in_rt_dat_data_d_1_118; // @[retiming.scala 9:92]
  reg [31:0] _RAND_118;
  reg [7:0] in_rt_dat_data_d_1_119; // @[retiming.scala 9:92]
  reg [31:0] _RAND_119;
  reg [7:0] in_rt_dat_data_d_1_120; // @[retiming.scala 9:92]
  reg [31:0] _RAND_120;
  reg [7:0] in_rt_dat_data_d_1_121; // @[retiming.scala 9:92]
  reg [31:0] _RAND_121;
  reg [7:0] in_rt_dat_data_d_1_122; // @[retiming.scala 9:92]
  reg [31:0] _RAND_122;
  reg [7:0] in_rt_dat_data_d_1_123; // @[retiming.scala 9:92]
  reg [31:0] _RAND_123;
  reg [7:0] in_rt_dat_data_d_1_124; // @[retiming.scala 9:92]
  reg [31:0] _RAND_124;
  reg [7:0] in_rt_dat_data_d_1_125; // @[retiming.scala 9:92]
  reg [31:0] _RAND_125;
  reg [7:0] in_rt_dat_data_d_1_126; // @[retiming.scala 9:92]
  reg [31:0] _RAND_126;
  reg [7:0] in_rt_dat_data_d_1_127; // @[retiming.scala 9:92]
  reg [31:0] _RAND_127;
  reg [7:0] in_rt_dat_data_d_2_0; // @[retiming.scala 9:92]
  reg [31:0] _RAND_128;
  reg [7:0] in_rt_dat_data_d_2_1; // @[retiming.scala 9:92]
  reg [31:0] _RAND_129;
  reg [7:0] in_rt_dat_data_d_2_2; // @[retiming.scala 9:92]
  reg [31:0] _RAND_130;
  reg [7:0] in_rt_dat_data_d_2_3; // @[retiming.scala 9:92]
  reg [31:0] _RAND_131;
  reg [7:0] in_rt_dat_data_d_2_4; // @[retiming.scala 9:92]
  reg [31:0] _RAND_132;
  reg [7:0] in_rt_dat_data_d_2_5; // @[retiming.scala 9:92]
  reg [31:0] _RAND_133;
  reg [7:0] in_rt_dat_data_d_2_6; // @[retiming.scala 9:92]
  reg [31:0] _RAND_134;
  reg [7:0] in_rt_dat_data_d_2_7; // @[retiming.scala 9:92]
  reg [31:0] _RAND_135;
  reg [7:0] in_rt_dat_data_d_2_8; // @[retiming.scala 9:92]
  reg [31:0] _RAND_136;
  reg [7:0] in_rt_dat_data_d_2_9; // @[retiming.scala 9:92]
  reg [31:0] _RAND_137;
  reg [7:0] in_rt_dat_data_d_2_10; // @[retiming.scala 9:92]
  reg [31:0] _RAND_138;
  reg [7:0] in_rt_dat_data_d_2_11; // @[retiming.scala 9:92]
  reg [31:0] _RAND_139;
  reg [7:0] in_rt_dat_data_d_2_12; // @[retiming.scala 9:92]
  reg [31:0] _RAND_140;
  reg [7:0] in_rt_dat_data_d_2_13; // @[retiming.scala 9:92]
  reg [31:0] _RAND_141;
  reg [7:0] in_rt_dat_data_d_2_14; // @[retiming.scala 9:92]
  reg [31:0] _RAND_142;
  reg [7:0] in_rt_dat_data_d_2_15; // @[retiming.scala 9:92]
  reg [31:0] _RAND_143;
  reg [7:0] in_rt_dat_data_d_2_16; // @[retiming.scala 9:92]
  reg [31:0] _RAND_144;
  reg [7:0] in_rt_dat_data_d_2_17; // @[retiming.scala 9:92]
  reg [31:0] _RAND_145;
  reg [7:0] in_rt_dat_data_d_2_18; // @[retiming.scala 9:92]
  reg [31:0] _RAND_146;
  reg [7:0] in_rt_dat_data_d_2_19; // @[retiming.scala 9:92]
  reg [31:0] _RAND_147;
  reg [7:0] in_rt_dat_data_d_2_20; // @[retiming.scala 9:92]
  reg [31:0] _RAND_148;
  reg [7:0] in_rt_dat_data_d_2_21; // @[retiming.scala 9:92]
  reg [31:0] _RAND_149;
  reg [7:0] in_rt_dat_data_d_2_22; // @[retiming.scala 9:92]
  reg [31:0] _RAND_150;
  reg [7:0] in_rt_dat_data_d_2_23; // @[retiming.scala 9:92]
  reg [31:0] _RAND_151;
  reg [7:0] in_rt_dat_data_d_2_24; // @[retiming.scala 9:92]
  reg [31:0] _RAND_152;
  reg [7:0] in_rt_dat_data_d_2_25; // @[retiming.scala 9:92]
  reg [31:0] _RAND_153;
  reg [7:0] in_rt_dat_data_d_2_26; // @[retiming.scala 9:92]
  reg [31:0] _RAND_154;
  reg [7:0] in_rt_dat_data_d_2_27; // @[retiming.scala 9:92]
  reg [31:0] _RAND_155;
  reg [7:0] in_rt_dat_data_d_2_28; // @[retiming.scala 9:92]
  reg [31:0] _RAND_156;
  reg [7:0] in_rt_dat_data_d_2_29; // @[retiming.scala 9:92]
  reg [31:0] _RAND_157;
  reg [7:0] in_rt_dat_data_d_2_30; // @[retiming.scala 9:92]
  reg [31:0] _RAND_158;
  reg [7:0] in_rt_dat_data_d_2_31; // @[retiming.scala 9:92]
  reg [31:0] _RAND_159;
  reg [7:0] in_rt_dat_data_d_2_32; // @[retiming.scala 9:92]
  reg [31:0] _RAND_160;
  reg [7:0] in_rt_dat_data_d_2_33; // @[retiming.scala 9:92]
  reg [31:0] _RAND_161;
  reg [7:0] in_rt_dat_data_d_2_34; // @[retiming.scala 9:92]
  reg [31:0] _RAND_162;
  reg [7:0] in_rt_dat_data_d_2_35; // @[retiming.scala 9:92]
  reg [31:0] _RAND_163;
  reg [7:0] in_rt_dat_data_d_2_36; // @[retiming.scala 9:92]
  reg [31:0] _RAND_164;
  reg [7:0] in_rt_dat_data_d_2_37; // @[retiming.scala 9:92]
  reg [31:0] _RAND_165;
  reg [7:0] in_rt_dat_data_d_2_38; // @[retiming.scala 9:92]
  reg [31:0] _RAND_166;
  reg [7:0] in_rt_dat_data_d_2_39; // @[retiming.scala 9:92]
  reg [31:0] _RAND_167;
  reg [7:0] in_rt_dat_data_d_2_40; // @[retiming.scala 9:92]
  reg [31:0] _RAND_168;
  reg [7:0] in_rt_dat_data_d_2_41; // @[retiming.scala 9:92]
  reg [31:0] _RAND_169;
  reg [7:0] in_rt_dat_data_d_2_42; // @[retiming.scala 9:92]
  reg [31:0] _RAND_170;
  reg [7:0] in_rt_dat_data_d_2_43; // @[retiming.scala 9:92]
  reg [31:0] _RAND_171;
  reg [7:0] in_rt_dat_data_d_2_44; // @[retiming.scala 9:92]
  reg [31:0] _RAND_172;
  reg [7:0] in_rt_dat_data_d_2_45; // @[retiming.scala 9:92]
  reg [31:0] _RAND_173;
  reg [7:0] in_rt_dat_data_d_2_46; // @[retiming.scala 9:92]
  reg [31:0] _RAND_174;
  reg [7:0] in_rt_dat_data_d_2_47; // @[retiming.scala 9:92]
  reg [31:0] _RAND_175;
  reg [7:0] in_rt_dat_data_d_2_48; // @[retiming.scala 9:92]
  reg [31:0] _RAND_176;
  reg [7:0] in_rt_dat_data_d_2_49; // @[retiming.scala 9:92]
  reg [31:0] _RAND_177;
  reg [7:0] in_rt_dat_data_d_2_50; // @[retiming.scala 9:92]
  reg [31:0] _RAND_178;
  reg [7:0] in_rt_dat_data_d_2_51; // @[retiming.scala 9:92]
  reg [31:0] _RAND_179;
  reg [7:0] in_rt_dat_data_d_2_52; // @[retiming.scala 9:92]
  reg [31:0] _RAND_180;
  reg [7:0] in_rt_dat_data_d_2_53; // @[retiming.scala 9:92]
  reg [31:0] _RAND_181;
  reg [7:0] in_rt_dat_data_d_2_54; // @[retiming.scala 9:92]
  reg [31:0] _RAND_182;
  reg [7:0] in_rt_dat_data_d_2_55; // @[retiming.scala 9:92]
  reg [31:0] _RAND_183;
  reg [7:0] in_rt_dat_data_d_2_56; // @[retiming.scala 9:92]
  reg [31:0] _RAND_184;
  reg [7:0] in_rt_dat_data_d_2_57; // @[retiming.scala 9:92]
  reg [31:0] _RAND_185;
  reg [7:0] in_rt_dat_data_d_2_58; // @[retiming.scala 9:92]
  reg [31:0] _RAND_186;
  reg [7:0] in_rt_dat_data_d_2_59; // @[retiming.scala 9:92]
  reg [31:0] _RAND_187;
  reg [7:0] in_rt_dat_data_d_2_60; // @[retiming.scala 9:92]
  reg [31:0] _RAND_188;
  reg [7:0] in_rt_dat_data_d_2_61; // @[retiming.scala 9:92]
  reg [31:0] _RAND_189;
  reg [7:0] in_rt_dat_data_d_2_62; // @[retiming.scala 9:92]
  reg [31:0] _RAND_190;
  reg [7:0] in_rt_dat_data_d_2_63; // @[retiming.scala 9:92]
  reg [31:0] _RAND_191;
  reg [7:0] in_rt_dat_data_d_2_64; // @[retiming.scala 9:92]
  reg [31:0] _RAND_192;
  reg [7:0] in_rt_dat_data_d_2_65; // @[retiming.scala 9:92]
  reg [31:0] _RAND_193;
  reg [7:0] in_rt_dat_data_d_2_66; // @[retiming.scala 9:92]
  reg [31:0] _RAND_194;
  reg [7:0] in_rt_dat_data_d_2_67; // @[retiming.scala 9:92]
  reg [31:0] _RAND_195;
  reg [7:0] in_rt_dat_data_d_2_68; // @[retiming.scala 9:92]
  reg [31:0] _RAND_196;
  reg [7:0] in_rt_dat_data_d_2_69; // @[retiming.scala 9:92]
  reg [31:0] _RAND_197;
  reg [7:0] in_rt_dat_data_d_2_70; // @[retiming.scala 9:92]
  reg [31:0] _RAND_198;
  reg [7:0] in_rt_dat_data_d_2_71; // @[retiming.scala 9:92]
  reg [31:0] _RAND_199;
  reg [7:0] in_rt_dat_data_d_2_72; // @[retiming.scala 9:92]
  reg [31:0] _RAND_200;
  reg [7:0] in_rt_dat_data_d_2_73; // @[retiming.scala 9:92]
  reg [31:0] _RAND_201;
  reg [7:0] in_rt_dat_data_d_2_74; // @[retiming.scala 9:92]
  reg [31:0] _RAND_202;
  reg [7:0] in_rt_dat_data_d_2_75; // @[retiming.scala 9:92]
  reg [31:0] _RAND_203;
  reg [7:0] in_rt_dat_data_d_2_76; // @[retiming.scala 9:92]
  reg [31:0] _RAND_204;
  reg [7:0] in_rt_dat_data_d_2_77; // @[retiming.scala 9:92]
  reg [31:0] _RAND_205;
  reg [7:0] in_rt_dat_data_d_2_78; // @[retiming.scala 9:92]
  reg [31:0] _RAND_206;
  reg [7:0] in_rt_dat_data_d_2_79; // @[retiming.scala 9:92]
  reg [31:0] _RAND_207;
  reg [7:0] in_rt_dat_data_d_2_80; // @[retiming.scala 9:92]
  reg [31:0] _RAND_208;
  reg [7:0] in_rt_dat_data_d_2_81; // @[retiming.scala 9:92]
  reg [31:0] _RAND_209;
  reg [7:0] in_rt_dat_data_d_2_82; // @[retiming.scala 9:92]
  reg [31:0] _RAND_210;
  reg [7:0] in_rt_dat_data_d_2_83; // @[retiming.scala 9:92]
  reg [31:0] _RAND_211;
  reg [7:0] in_rt_dat_data_d_2_84; // @[retiming.scala 9:92]
  reg [31:0] _RAND_212;
  reg [7:0] in_rt_dat_data_d_2_85; // @[retiming.scala 9:92]
  reg [31:0] _RAND_213;
  reg [7:0] in_rt_dat_data_d_2_86; // @[retiming.scala 9:92]
  reg [31:0] _RAND_214;
  reg [7:0] in_rt_dat_data_d_2_87; // @[retiming.scala 9:92]
  reg [31:0] _RAND_215;
  reg [7:0] in_rt_dat_data_d_2_88; // @[retiming.scala 9:92]
  reg [31:0] _RAND_216;
  reg [7:0] in_rt_dat_data_d_2_89; // @[retiming.scala 9:92]
  reg [31:0] _RAND_217;
  reg [7:0] in_rt_dat_data_d_2_90; // @[retiming.scala 9:92]
  reg [31:0] _RAND_218;
  reg [7:0] in_rt_dat_data_d_2_91; // @[retiming.scala 9:92]
  reg [31:0] _RAND_219;
  reg [7:0] in_rt_dat_data_d_2_92; // @[retiming.scala 9:92]
  reg [31:0] _RAND_220;
  reg [7:0] in_rt_dat_data_d_2_93; // @[retiming.scala 9:92]
  reg [31:0] _RAND_221;
  reg [7:0] in_rt_dat_data_d_2_94; // @[retiming.scala 9:92]
  reg [31:0] _RAND_222;
  reg [7:0] in_rt_dat_data_d_2_95; // @[retiming.scala 9:92]
  reg [31:0] _RAND_223;
  reg [7:0] in_rt_dat_data_d_2_96; // @[retiming.scala 9:92]
  reg [31:0] _RAND_224;
  reg [7:0] in_rt_dat_data_d_2_97; // @[retiming.scala 9:92]
  reg [31:0] _RAND_225;
  reg [7:0] in_rt_dat_data_d_2_98; // @[retiming.scala 9:92]
  reg [31:0] _RAND_226;
  reg [7:0] in_rt_dat_data_d_2_99; // @[retiming.scala 9:92]
  reg [31:0] _RAND_227;
  reg [7:0] in_rt_dat_data_d_2_100; // @[retiming.scala 9:92]
  reg [31:0] _RAND_228;
  reg [7:0] in_rt_dat_data_d_2_101; // @[retiming.scala 9:92]
  reg [31:0] _RAND_229;
  reg [7:0] in_rt_dat_data_d_2_102; // @[retiming.scala 9:92]
  reg [31:0] _RAND_230;
  reg [7:0] in_rt_dat_data_d_2_103; // @[retiming.scala 9:92]
  reg [31:0] _RAND_231;
  reg [7:0] in_rt_dat_data_d_2_104; // @[retiming.scala 9:92]
  reg [31:0] _RAND_232;
  reg [7:0] in_rt_dat_data_d_2_105; // @[retiming.scala 9:92]
  reg [31:0] _RAND_233;
  reg [7:0] in_rt_dat_data_d_2_106; // @[retiming.scala 9:92]
  reg [31:0] _RAND_234;
  reg [7:0] in_rt_dat_data_d_2_107; // @[retiming.scala 9:92]
  reg [31:0] _RAND_235;
  reg [7:0] in_rt_dat_data_d_2_108; // @[retiming.scala 9:92]
  reg [31:0] _RAND_236;
  reg [7:0] in_rt_dat_data_d_2_109; // @[retiming.scala 9:92]
  reg [31:0] _RAND_237;
  reg [7:0] in_rt_dat_data_d_2_110; // @[retiming.scala 9:92]
  reg [31:0] _RAND_238;
  reg [7:0] in_rt_dat_data_d_2_111; // @[retiming.scala 9:92]
  reg [31:0] _RAND_239;
  reg [7:0] in_rt_dat_data_d_2_112; // @[retiming.scala 9:92]
  reg [31:0] _RAND_240;
  reg [7:0] in_rt_dat_data_d_2_113; // @[retiming.scala 9:92]
  reg [31:0] _RAND_241;
  reg [7:0] in_rt_dat_data_d_2_114; // @[retiming.scala 9:92]
  reg [31:0] _RAND_242;
  reg [7:0] in_rt_dat_data_d_2_115; // @[retiming.scala 9:92]
  reg [31:0] _RAND_243;
  reg [7:0] in_rt_dat_data_d_2_116; // @[retiming.scala 9:92]
  reg [31:0] _RAND_244;
  reg [7:0] in_rt_dat_data_d_2_117; // @[retiming.scala 9:92]
  reg [31:0] _RAND_245;
  reg [7:0] in_rt_dat_data_d_2_118; // @[retiming.scala 9:92]
  reg [31:0] _RAND_246;
  reg [7:0] in_rt_dat_data_d_2_119; // @[retiming.scala 9:92]
  reg [31:0] _RAND_247;
  reg [7:0] in_rt_dat_data_d_2_120; // @[retiming.scala 9:92]
  reg [31:0] _RAND_248;
  reg [7:0] in_rt_dat_data_d_2_121; // @[retiming.scala 9:92]
  reg [31:0] _RAND_249;
  reg [7:0] in_rt_dat_data_d_2_122; // @[retiming.scala 9:92]
  reg [31:0] _RAND_250;
  reg [7:0] in_rt_dat_data_d_2_123; // @[retiming.scala 9:92]
  reg [31:0] _RAND_251;
  reg [7:0] in_rt_dat_data_d_2_124; // @[retiming.scala 9:92]
  reg [31:0] _RAND_252;
  reg [7:0] in_rt_dat_data_d_2_125; // @[retiming.scala 9:92]
  reg [31:0] _RAND_253;
  reg [7:0] in_rt_dat_data_d_2_126; // @[retiming.scala 9:92]
  reg [31:0] _RAND_254;
  reg [7:0] in_rt_dat_data_d_2_127; // @[retiming.scala 9:92]
  reg [31:0] _RAND_255;
  reg  in_rt_dat_mask_d_1_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_256;
  reg  in_rt_dat_mask_d_1_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_257;
  reg  in_rt_dat_mask_d_1_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_258;
  reg  in_rt_dat_mask_d_1_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_259;
  reg  in_rt_dat_mask_d_1_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_260;
  reg  in_rt_dat_mask_d_1_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_261;
  reg  in_rt_dat_mask_d_1_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_262;
  reg  in_rt_dat_mask_d_1_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_263;
  reg  in_rt_dat_mask_d_1_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_264;
  reg  in_rt_dat_mask_d_1_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_265;
  reg  in_rt_dat_mask_d_1_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_266;
  reg  in_rt_dat_mask_d_1_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_267;
  reg  in_rt_dat_mask_d_1_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_268;
  reg  in_rt_dat_mask_d_1_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_269;
  reg  in_rt_dat_mask_d_1_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_270;
  reg  in_rt_dat_mask_d_1_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_271;
  reg  in_rt_dat_mask_d_1_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_272;
  reg  in_rt_dat_mask_d_1_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_273;
  reg  in_rt_dat_mask_d_1_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_274;
  reg  in_rt_dat_mask_d_1_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_275;
  reg  in_rt_dat_mask_d_1_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_276;
  reg  in_rt_dat_mask_d_1_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_277;
  reg  in_rt_dat_mask_d_1_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_278;
  reg  in_rt_dat_mask_d_1_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_279;
  reg  in_rt_dat_mask_d_1_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_280;
  reg  in_rt_dat_mask_d_1_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_281;
  reg  in_rt_dat_mask_d_1_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_282;
  reg  in_rt_dat_mask_d_1_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_283;
  reg  in_rt_dat_mask_d_1_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_284;
  reg  in_rt_dat_mask_d_1_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_285;
  reg  in_rt_dat_mask_d_1_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_286;
  reg  in_rt_dat_mask_d_1_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_287;
  reg  in_rt_dat_mask_d_1_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_288;
  reg  in_rt_dat_mask_d_1_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_289;
  reg  in_rt_dat_mask_d_1_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_290;
  reg  in_rt_dat_mask_d_1_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_291;
  reg  in_rt_dat_mask_d_1_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_292;
  reg  in_rt_dat_mask_d_1_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_293;
  reg  in_rt_dat_mask_d_1_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_294;
  reg  in_rt_dat_mask_d_1_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_295;
  reg  in_rt_dat_mask_d_1_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_296;
  reg  in_rt_dat_mask_d_1_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_297;
  reg  in_rt_dat_mask_d_1_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_298;
  reg  in_rt_dat_mask_d_1_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_299;
  reg  in_rt_dat_mask_d_1_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_300;
  reg  in_rt_dat_mask_d_1_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_301;
  reg  in_rt_dat_mask_d_1_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_302;
  reg  in_rt_dat_mask_d_1_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_303;
  reg  in_rt_dat_mask_d_1_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_304;
  reg  in_rt_dat_mask_d_1_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_305;
  reg  in_rt_dat_mask_d_1_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_306;
  reg  in_rt_dat_mask_d_1_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_307;
  reg  in_rt_dat_mask_d_1_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_308;
  reg  in_rt_dat_mask_d_1_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_309;
  reg  in_rt_dat_mask_d_1_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_310;
  reg  in_rt_dat_mask_d_1_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_311;
  reg  in_rt_dat_mask_d_1_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_312;
  reg  in_rt_dat_mask_d_1_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_313;
  reg  in_rt_dat_mask_d_1_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_314;
  reg  in_rt_dat_mask_d_1_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_315;
  reg  in_rt_dat_mask_d_1_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_316;
  reg  in_rt_dat_mask_d_1_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_317;
  reg  in_rt_dat_mask_d_1_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_318;
  reg  in_rt_dat_mask_d_1_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_319;
  reg  in_rt_dat_mask_d_1_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_320;
  reg  in_rt_dat_mask_d_1_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_321;
  reg  in_rt_dat_mask_d_1_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_322;
  reg  in_rt_dat_mask_d_1_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_323;
  reg  in_rt_dat_mask_d_1_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_324;
  reg  in_rt_dat_mask_d_1_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_325;
  reg  in_rt_dat_mask_d_1_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_326;
  reg  in_rt_dat_mask_d_1_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_327;
  reg  in_rt_dat_mask_d_1_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_328;
  reg  in_rt_dat_mask_d_1_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_329;
  reg  in_rt_dat_mask_d_1_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_330;
  reg  in_rt_dat_mask_d_1_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_331;
  reg  in_rt_dat_mask_d_1_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_332;
  reg  in_rt_dat_mask_d_1_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_333;
  reg  in_rt_dat_mask_d_1_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_334;
  reg  in_rt_dat_mask_d_1_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_335;
  reg  in_rt_dat_mask_d_1_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_336;
  reg  in_rt_dat_mask_d_1_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_337;
  reg  in_rt_dat_mask_d_1_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_338;
  reg  in_rt_dat_mask_d_1_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_339;
  reg  in_rt_dat_mask_d_1_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_340;
  reg  in_rt_dat_mask_d_1_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_341;
  reg  in_rt_dat_mask_d_1_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_342;
  reg  in_rt_dat_mask_d_1_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_343;
  reg  in_rt_dat_mask_d_1_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_344;
  reg  in_rt_dat_mask_d_1_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_345;
  reg  in_rt_dat_mask_d_1_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_346;
  reg  in_rt_dat_mask_d_1_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_347;
  reg  in_rt_dat_mask_d_1_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_348;
  reg  in_rt_dat_mask_d_1_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_349;
  reg  in_rt_dat_mask_d_1_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_350;
  reg  in_rt_dat_mask_d_1_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_351;
  reg  in_rt_dat_mask_d_1_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_352;
  reg  in_rt_dat_mask_d_1_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_353;
  reg  in_rt_dat_mask_d_1_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_354;
  reg  in_rt_dat_mask_d_1_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_355;
  reg  in_rt_dat_mask_d_1_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_356;
  reg  in_rt_dat_mask_d_1_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_357;
  reg  in_rt_dat_mask_d_1_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_358;
  reg  in_rt_dat_mask_d_1_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_359;
  reg  in_rt_dat_mask_d_1_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_360;
  reg  in_rt_dat_mask_d_1_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_361;
  reg  in_rt_dat_mask_d_1_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_362;
  reg  in_rt_dat_mask_d_1_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_363;
  reg  in_rt_dat_mask_d_1_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_364;
  reg  in_rt_dat_mask_d_1_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_365;
  reg  in_rt_dat_mask_d_1_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_366;
  reg  in_rt_dat_mask_d_1_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_367;
  reg  in_rt_dat_mask_d_1_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_368;
  reg  in_rt_dat_mask_d_1_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_369;
  reg  in_rt_dat_mask_d_1_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_370;
  reg  in_rt_dat_mask_d_1_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_371;
  reg  in_rt_dat_mask_d_1_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_372;
  reg  in_rt_dat_mask_d_1_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_373;
  reg  in_rt_dat_mask_d_1_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_374;
  reg  in_rt_dat_mask_d_1_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_375;
  reg  in_rt_dat_mask_d_1_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_376;
  reg  in_rt_dat_mask_d_1_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_377;
  reg  in_rt_dat_mask_d_1_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_378;
  reg  in_rt_dat_mask_d_1_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_379;
  reg  in_rt_dat_mask_d_1_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_380;
  reg  in_rt_dat_mask_d_1_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_381;
  reg  in_rt_dat_mask_d_1_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_382;
  reg  in_rt_dat_mask_d_1_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_383;
  reg  in_rt_dat_mask_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_384;
  reg  in_rt_dat_mask_d_2_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_385;
  reg  in_rt_dat_mask_d_2_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_386;
  reg  in_rt_dat_mask_d_2_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_387;
  reg  in_rt_dat_mask_d_2_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_388;
  reg  in_rt_dat_mask_d_2_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_389;
  reg  in_rt_dat_mask_d_2_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_390;
  reg  in_rt_dat_mask_d_2_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_391;
  reg  in_rt_dat_mask_d_2_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_392;
  reg  in_rt_dat_mask_d_2_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_393;
  reg  in_rt_dat_mask_d_2_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_394;
  reg  in_rt_dat_mask_d_2_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_395;
  reg  in_rt_dat_mask_d_2_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_396;
  reg  in_rt_dat_mask_d_2_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_397;
  reg  in_rt_dat_mask_d_2_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_398;
  reg  in_rt_dat_mask_d_2_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_399;
  reg  in_rt_dat_mask_d_2_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_400;
  reg  in_rt_dat_mask_d_2_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_401;
  reg  in_rt_dat_mask_d_2_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_402;
  reg  in_rt_dat_mask_d_2_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_403;
  reg  in_rt_dat_mask_d_2_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_404;
  reg  in_rt_dat_mask_d_2_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_405;
  reg  in_rt_dat_mask_d_2_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_406;
  reg  in_rt_dat_mask_d_2_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_407;
  reg  in_rt_dat_mask_d_2_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_408;
  reg  in_rt_dat_mask_d_2_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_409;
  reg  in_rt_dat_mask_d_2_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_410;
  reg  in_rt_dat_mask_d_2_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_411;
  reg  in_rt_dat_mask_d_2_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_412;
  reg  in_rt_dat_mask_d_2_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_413;
  reg  in_rt_dat_mask_d_2_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_414;
  reg  in_rt_dat_mask_d_2_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_415;
  reg  in_rt_dat_mask_d_2_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_416;
  reg  in_rt_dat_mask_d_2_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_417;
  reg  in_rt_dat_mask_d_2_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_418;
  reg  in_rt_dat_mask_d_2_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_419;
  reg  in_rt_dat_mask_d_2_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_420;
  reg  in_rt_dat_mask_d_2_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_421;
  reg  in_rt_dat_mask_d_2_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_422;
  reg  in_rt_dat_mask_d_2_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_423;
  reg  in_rt_dat_mask_d_2_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_424;
  reg  in_rt_dat_mask_d_2_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_425;
  reg  in_rt_dat_mask_d_2_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_426;
  reg  in_rt_dat_mask_d_2_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_427;
  reg  in_rt_dat_mask_d_2_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_428;
  reg  in_rt_dat_mask_d_2_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_429;
  reg  in_rt_dat_mask_d_2_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_430;
  reg  in_rt_dat_mask_d_2_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_431;
  reg  in_rt_dat_mask_d_2_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_432;
  reg  in_rt_dat_mask_d_2_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_433;
  reg  in_rt_dat_mask_d_2_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_434;
  reg  in_rt_dat_mask_d_2_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_435;
  reg  in_rt_dat_mask_d_2_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_436;
  reg  in_rt_dat_mask_d_2_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_437;
  reg  in_rt_dat_mask_d_2_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_438;
  reg  in_rt_dat_mask_d_2_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_439;
  reg  in_rt_dat_mask_d_2_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_440;
  reg  in_rt_dat_mask_d_2_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_441;
  reg  in_rt_dat_mask_d_2_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_442;
  reg  in_rt_dat_mask_d_2_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_443;
  reg  in_rt_dat_mask_d_2_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_444;
  reg  in_rt_dat_mask_d_2_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_445;
  reg  in_rt_dat_mask_d_2_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_446;
  reg  in_rt_dat_mask_d_2_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_447;
  reg  in_rt_dat_mask_d_2_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_448;
  reg  in_rt_dat_mask_d_2_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_449;
  reg  in_rt_dat_mask_d_2_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_450;
  reg  in_rt_dat_mask_d_2_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_451;
  reg  in_rt_dat_mask_d_2_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_452;
  reg  in_rt_dat_mask_d_2_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_453;
  reg  in_rt_dat_mask_d_2_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_454;
  reg  in_rt_dat_mask_d_2_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_455;
  reg  in_rt_dat_mask_d_2_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_456;
  reg  in_rt_dat_mask_d_2_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_457;
  reg  in_rt_dat_mask_d_2_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_458;
  reg  in_rt_dat_mask_d_2_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_459;
  reg  in_rt_dat_mask_d_2_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_460;
  reg  in_rt_dat_mask_d_2_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_461;
  reg  in_rt_dat_mask_d_2_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_462;
  reg  in_rt_dat_mask_d_2_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_463;
  reg  in_rt_dat_mask_d_2_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_464;
  reg  in_rt_dat_mask_d_2_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_465;
  reg  in_rt_dat_mask_d_2_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_466;
  reg  in_rt_dat_mask_d_2_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_467;
  reg  in_rt_dat_mask_d_2_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_468;
  reg  in_rt_dat_mask_d_2_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_469;
  reg  in_rt_dat_mask_d_2_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_470;
  reg  in_rt_dat_mask_d_2_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_471;
  reg  in_rt_dat_mask_d_2_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_472;
  reg  in_rt_dat_mask_d_2_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_473;
  reg  in_rt_dat_mask_d_2_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_474;
  reg  in_rt_dat_mask_d_2_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_475;
  reg  in_rt_dat_mask_d_2_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_476;
  reg  in_rt_dat_mask_d_2_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_477;
  reg  in_rt_dat_mask_d_2_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_478;
  reg  in_rt_dat_mask_d_2_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_479;
  reg  in_rt_dat_mask_d_2_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_480;
  reg  in_rt_dat_mask_d_2_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_481;
  reg  in_rt_dat_mask_d_2_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_482;
  reg  in_rt_dat_mask_d_2_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_483;
  reg  in_rt_dat_mask_d_2_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_484;
  reg  in_rt_dat_mask_d_2_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_485;
  reg  in_rt_dat_mask_d_2_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_486;
  reg  in_rt_dat_mask_d_2_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_487;
  reg  in_rt_dat_mask_d_2_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_488;
  reg  in_rt_dat_mask_d_2_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_489;
  reg  in_rt_dat_mask_d_2_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_490;
  reg  in_rt_dat_mask_d_2_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_491;
  reg  in_rt_dat_mask_d_2_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_492;
  reg  in_rt_dat_mask_d_2_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_493;
  reg  in_rt_dat_mask_d_2_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_494;
  reg  in_rt_dat_mask_d_2_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_495;
  reg  in_rt_dat_mask_d_2_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_496;
  reg  in_rt_dat_mask_d_2_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_497;
  reg  in_rt_dat_mask_d_2_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_498;
  reg  in_rt_dat_mask_d_2_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_499;
  reg  in_rt_dat_mask_d_2_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_500;
  reg  in_rt_dat_mask_d_2_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_501;
  reg  in_rt_dat_mask_d_2_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_502;
  reg  in_rt_dat_mask_d_2_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_503;
  reg  in_rt_dat_mask_d_2_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_504;
  reg  in_rt_dat_mask_d_2_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_505;
  reg  in_rt_dat_mask_d_2_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_506;
  reg  in_rt_dat_mask_d_2_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_507;
  reg  in_rt_dat_mask_d_2_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_508;
  reg  in_rt_dat_mask_d_2_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_509;
  reg  in_rt_dat_mask_d_2_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_510;
  reg  in_rt_dat_mask_d_2_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 60:70]
  reg [31:0] _RAND_511;
  reg  in_rt_dat_pvld_d_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 62:70]
  reg [31:0] _RAND_512;
  reg  in_rt_dat_pvld_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 62:70]
  reg [31:0] _RAND_513;
  reg [8:0] in_rt_dat_pd_d_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 64:70]
  reg [31:0] _RAND_514;
  reg [8:0] in_rt_dat_pd_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 64:70]
  reg [31:0] _RAND_515;
  reg [7:0] in_rt_wt_data_d_1_0; // @[retiming.scala 9:92]
  reg [31:0] _RAND_516;
  reg [7:0] in_rt_wt_data_d_1_1; // @[retiming.scala 9:92]
  reg [31:0] _RAND_517;
  reg [7:0] in_rt_wt_data_d_1_2; // @[retiming.scala 9:92]
  reg [31:0] _RAND_518;
  reg [7:0] in_rt_wt_data_d_1_3; // @[retiming.scala 9:92]
  reg [31:0] _RAND_519;
  reg [7:0] in_rt_wt_data_d_1_4; // @[retiming.scala 9:92]
  reg [31:0] _RAND_520;
  reg [7:0] in_rt_wt_data_d_1_5; // @[retiming.scala 9:92]
  reg [31:0] _RAND_521;
  reg [7:0] in_rt_wt_data_d_1_6; // @[retiming.scala 9:92]
  reg [31:0] _RAND_522;
  reg [7:0] in_rt_wt_data_d_1_7; // @[retiming.scala 9:92]
  reg [31:0] _RAND_523;
  reg [7:0] in_rt_wt_data_d_1_8; // @[retiming.scala 9:92]
  reg [31:0] _RAND_524;
  reg [7:0] in_rt_wt_data_d_1_9; // @[retiming.scala 9:92]
  reg [31:0] _RAND_525;
  reg [7:0] in_rt_wt_data_d_1_10; // @[retiming.scala 9:92]
  reg [31:0] _RAND_526;
  reg [7:0] in_rt_wt_data_d_1_11; // @[retiming.scala 9:92]
  reg [31:0] _RAND_527;
  reg [7:0] in_rt_wt_data_d_1_12; // @[retiming.scala 9:92]
  reg [31:0] _RAND_528;
  reg [7:0] in_rt_wt_data_d_1_13; // @[retiming.scala 9:92]
  reg [31:0] _RAND_529;
  reg [7:0] in_rt_wt_data_d_1_14; // @[retiming.scala 9:92]
  reg [31:0] _RAND_530;
  reg [7:0] in_rt_wt_data_d_1_15; // @[retiming.scala 9:92]
  reg [31:0] _RAND_531;
  reg [7:0] in_rt_wt_data_d_1_16; // @[retiming.scala 9:92]
  reg [31:0] _RAND_532;
  reg [7:0] in_rt_wt_data_d_1_17; // @[retiming.scala 9:92]
  reg [31:0] _RAND_533;
  reg [7:0] in_rt_wt_data_d_1_18; // @[retiming.scala 9:92]
  reg [31:0] _RAND_534;
  reg [7:0] in_rt_wt_data_d_1_19; // @[retiming.scala 9:92]
  reg [31:0] _RAND_535;
  reg [7:0] in_rt_wt_data_d_1_20; // @[retiming.scala 9:92]
  reg [31:0] _RAND_536;
  reg [7:0] in_rt_wt_data_d_1_21; // @[retiming.scala 9:92]
  reg [31:0] _RAND_537;
  reg [7:0] in_rt_wt_data_d_1_22; // @[retiming.scala 9:92]
  reg [31:0] _RAND_538;
  reg [7:0] in_rt_wt_data_d_1_23; // @[retiming.scala 9:92]
  reg [31:0] _RAND_539;
  reg [7:0] in_rt_wt_data_d_1_24; // @[retiming.scala 9:92]
  reg [31:0] _RAND_540;
  reg [7:0] in_rt_wt_data_d_1_25; // @[retiming.scala 9:92]
  reg [31:0] _RAND_541;
  reg [7:0] in_rt_wt_data_d_1_26; // @[retiming.scala 9:92]
  reg [31:0] _RAND_542;
  reg [7:0] in_rt_wt_data_d_1_27; // @[retiming.scala 9:92]
  reg [31:0] _RAND_543;
  reg [7:0] in_rt_wt_data_d_1_28; // @[retiming.scala 9:92]
  reg [31:0] _RAND_544;
  reg [7:0] in_rt_wt_data_d_1_29; // @[retiming.scala 9:92]
  reg [31:0] _RAND_545;
  reg [7:0] in_rt_wt_data_d_1_30; // @[retiming.scala 9:92]
  reg [31:0] _RAND_546;
  reg [7:0] in_rt_wt_data_d_1_31; // @[retiming.scala 9:92]
  reg [31:0] _RAND_547;
  reg [7:0] in_rt_wt_data_d_1_32; // @[retiming.scala 9:92]
  reg [31:0] _RAND_548;
  reg [7:0] in_rt_wt_data_d_1_33; // @[retiming.scala 9:92]
  reg [31:0] _RAND_549;
  reg [7:0] in_rt_wt_data_d_1_34; // @[retiming.scala 9:92]
  reg [31:0] _RAND_550;
  reg [7:0] in_rt_wt_data_d_1_35; // @[retiming.scala 9:92]
  reg [31:0] _RAND_551;
  reg [7:0] in_rt_wt_data_d_1_36; // @[retiming.scala 9:92]
  reg [31:0] _RAND_552;
  reg [7:0] in_rt_wt_data_d_1_37; // @[retiming.scala 9:92]
  reg [31:0] _RAND_553;
  reg [7:0] in_rt_wt_data_d_1_38; // @[retiming.scala 9:92]
  reg [31:0] _RAND_554;
  reg [7:0] in_rt_wt_data_d_1_39; // @[retiming.scala 9:92]
  reg [31:0] _RAND_555;
  reg [7:0] in_rt_wt_data_d_1_40; // @[retiming.scala 9:92]
  reg [31:0] _RAND_556;
  reg [7:0] in_rt_wt_data_d_1_41; // @[retiming.scala 9:92]
  reg [31:0] _RAND_557;
  reg [7:0] in_rt_wt_data_d_1_42; // @[retiming.scala 9:92]
  reg [31:0] _RAND_558;
  reg [7:0] in_rt_wt_data_d_1_43; // @[retiming.scala 9:92]
  reg [31:0] _RAND_559;
  reg [7:0] in_rt_wt_data_d_1_44; // @[retiming.scala 9:92]
  reg [31:0] _RAND_560;
  reg [7:0] in_rt_wt_data_d_1_45; // @[retiming.scala 9:92]
  reg [31:0] _RAND_561;
  reg [7:0] in_rt_wt_data_d_1_46; // @[retiming.scala 9:92]
  reg [31:0] _RAND_562;
  reg [7:0] in_rt_wt_data_d_1_47; // @[retiming.scala 9:92]
  reg [31:0] _RAND_563;
  reg [7:0] in_rt_wt_data_d_1_48; // @[retiming.scala 9:92]
  reg [31:0] _RAND_564;
  reg [7:0] in_rt_wt_data_d_1_49; // @[retiming.scala 9:92]
  reg [31:0] _RAND_565;
  reg [7:0] in_rt_wt_data_d_1_50; // @[retiming.scala 9:92]
  reg [31:0] _RAND_566;
  reg [7:0] in_rt_wt_data_d_1_51; // @[retiming.scala 9:92]
  reg [31:0] _RAND_567;
  reg [7:0] in_rt_wt_data_d_1_52; // @[retiming.scala 9:92]
  reg [31:0] _RAND_568;
  reg [7:0] in_rt_wt_data_d_1_53; // @[retiming.scala 9:92]
  reg [31:0] _RAND_569;
  reg [7:0] in_rt_wt_data_d_1_54; // @[retiming.scala 9:92]
  reg [31:0] _RAND_570;
  reg [7:0] in_rt_wt_data_d_1_55; // @[retiming.scala 9:92]
  reg [31:0] _RAND_571;
  reg [7:0] in_rt_wt_data_d_1_56; // @[retiming.scala 9:92]
  reg [31:0] _RAND_572;
  reg [7:0] in_rt_wt_data_d_1_57; // @[retiming.scala 9:92]
  reg [31:0] _RAND_573;
  reg [7:0] in_rt_wt_data_d_1_58; // @[retiming.scala 9:92]
  reg [31:0] _RAND_574;
  reg [7:0] in_rt_wt_data_d_1_59; // @[retiming.scala 9:92]
  reg [31:0] _RAND_575;
  reg [7:0] in_rt_wt_data_d_1_60; // @[retiming.scala 9:92]
  reg [31:0] _RAND_576;
  reg [7:0] in_rt_wt_data_d_1_61; // @[retiming.scala 9:92]
  reg [31:0] _RAND_577;
  reg [7:0] in_rt_wt_data_d_1_62; // @[retiming.scala 9:92]
  reg [31:0] _RAND_578;
  reg [7:0] in_rt_wt_data_d_1_63; // @[retiming.scala 9:92]
  reg [31:0] _RAND_579;
  reg [7:0] in_rt_wt_data_d_1_64; // @[retiming.scala 9:92]
  reg [31:0] _RAND_580;
  reg [7:0] in_rt_wt_data_d_1_65; // @[retiming.scala 9:92]
  reg [31:0] _RAND_581;
  reg [7:0] in_rt_wt_data_d_1_66; // @[retiming.scala 9:92]
  reg [31:0] _RAND_582;
  reg [7:0] in_rt_wt_data_d_1_67; // @[retiming.scala 9:92]
  reg [31:0] _RAND_583;
  reg [7:0] in_rt_wt_data_d_1_68; // @[retiming.scala 9:92]
  reg [31:0] _RAND_584;
  reg [7:0] in_rt_wt_data_d_1_69; // @[retiming.scala 9:92]
  reg [31:0] _RAND_585;
  reg [7:0] in_rt_wt_data_d_1_70; // @[retiming.scala 9:92]
  reg [31:0] _RAND_586;
  reg [7:0] in_rt_wt_data_d_1_71; // @[retiming.scala 9:92]
  reg [31:0] _RAND_587;
  reg [7:0] in_rt_wt_data_d_1_72; // @[retiming.scala 9:92]
  reg [31:0] _RAND_588;
  reg [7:0] in_rt_wt_data_d_1_73; // @[retiming.scala 9:92]
  reg [31:0] _RAND_589;
  reg [7:0] in_rt_wt_data_d_1_74; // @[retiming.scala 9:92]
  reg [31:0] _RAND_590;
  reg [7:0] in_rt_wt_data_d_1_75; // @[retiming.scala 9:92]
  reg [31:0] _RAND_591;
  reg [7:0] in_rt_wt_data_d_1_76; // @[retiming.scala 9:92]
  reg [31:0] _RAND_592;
  reg [7:0] in_rt_wt_data_d_1_77; // @[retiming.scala 9:92]
  reg [31:0] _RAND_593;
  reg [7:0] in_rt_wt_data_d_1_78; // @[retiming.scala 9:92]
  reg [31:0] _RAND_594;
  reg [7:0] in_rt_wt_data_d_1_79; // @[retiming.scala 9:92]
  reg [31:0] _RAND_595;
  reg [7:0] in_rt_wt_data_d_1_80; // @[retiming.scala 9:92]
  reg [31:0] _RAND_596;
  reg [7:0] in_rt_wt_data_d_1_81; // @[retiming.scala 9:92]
  reg [31:0] _RAND_597;
  reg [7:0] in_rt_wt_data_d_1_82; // @[retiming.scala 9:92]
  reg [31:0] _RAND_598;
  reg [7:0] in_rt_wt_data_d_1_83; // @[retiming.scala 9:92]
  reg [31:0] _RAND_599;
  reg [7:0] in_rt_wt_data_d_1_84; // @[retiming.scala 9:92]
  reg [31:0] _RAND_600;
  reg [7:0] in_rt_wt_data_d_1_85; // @[retiming.scala 9:92]
  reg [31:0] _RAND_601;
  reg [7:0] in_rt_wt_data_d_1_86; // @[retiming.scala 9:92]
  reg [31:0] _RAND_602;
  reg [7:0] in_rt_wt_data_d_1_87; // @[retiming.scala 9:92]
  reg [31:0] _RAND_603;
  reg [7:0] in_rt_wt_data_d_1_88; // @[retiming.scala 9:92]
  reg [31:0] _RAND_604;
  reg [7:0] in_rt_wt_data_d_1_89; // @[retiming.scala 9:92]
  reg [31:0] _RAND_605;
  reg [7:0] in_rt_wt_data_d_1_90; // @[retiming.scala 9:92]
  reg [31:0] _RAND_606;
  reg [7:0] in_rt_wt_data_d_1_91; // @[retiming.scala 9:92]
  reg [31:0] _RAND_607;
  reg [7:0] in_rt_wt_data_d_1_92; // @[retiming.scala 9:92]
  reg [31:0] _RAND_608;
  reg [7:0] in_rt_wt_data_d_1_93; // @[retiming.scala 9:92]
  reg [31:0] _RAND_609;
  reg [7:0] in_rt_wt_data_d_1_94; // @[retiming.scala 9:92]
  reg [31:0] _RAND_610;
  reg [7:0] in_rt_wt_data_d_1_95; // @[retiming.scala 9:92]
  reg [31:0] _RAND_611;
  reg [7:0] in_rt_wt_data_d_1_96; // @[retiming.scala 9:92]
  reg [31:0] _RAND_612;
  reg [7:0] in_rt_wt_data_d_1_97; // @[retiming.scala 9:92]
  reg [31:0] _RAND_613;
  reg [7:0] in_rt_wt_data_d_1_98; // @[retiming.scala 9:92]
  reg [31:0] _RAND_614;
  reg [7:0] in_rt_wt_data_d_1_99; // @[retiming.scala 9:92]
  reg [31:0] _RAND_615;
  reg [7:0] in_rt_wt_data_d_1_100; // @[retiming.scala 9:92]
  reg [31:0] _RAND_616;
  reg [7:0] in_rt_wt_data_d_1_101; // @[retiming.scala 9:92]
  reg [31:0] _RAND_617;
  reg [7:0] in_rt_wt_data_d_1_102; // @[retiming.scala 9:92]
  reg [31:0] _RAND_618;
  reg [7:0] in_rt_wt_data_d_1_103; // @[retiming.scala 9:92]
  reg [31:0] _RAND_619;
  reg [7:0] in_rt_wt_data_d_1_104; // @[retiming.scala 9:92]
  reg [31:0] _RAND_620;
  reg [7:0] in_rt_wt_data_d_1_105; // @[retiming.scala 9:92]
  reg [31:0] _RAND_621;
  reg [7:0] in_rt_wt_data_d_1_106; // @[retiming.scala 9:92]
  reg [31:0] _RAND_622;
  reg [7:0] in_rt_wt_data_d_1_107; // @[retiming.scala 9:92]
  reg [31:0] _RAND_623;
  reg [7:0] in_rt_wt_data_d_1_108; // @[retiming.scala 9:92]
  reg [31:0] _RAND_624;
  reg [7:0] in_rt_wt_data_d_1_109; // @[retiming.scala 9:92]
  reg [31:0] _RAND_625;
  reg [7:0] in_rt_wt_data_d_1_110; // @[retiming.scala 9:92]
  reg [31:0] _RAND_626;
  reg [7:0] in_rt_wt_data_d_1_111; // @[retiming.scala 9:92]
  reg [31:0] _RAND_627;
  reg [7:0] in_rt_wt_data_d_1_112; // @[retiming.scala 9:92]
  reg [31:0] _RAND_628;
  reg [7:0] in_rt_wt_data_d_1_113; // @[retiming.scala 9:92]
  reg [31:0] _RAND_629;
  reg [7:0] in_rt_wt_data_d_1_114; // @[retiming.scala 9:92]
  reg [31:0] _RAND_630;
  reg [7:0] in_rt_wt_data_d_1_115; // @[retiming.scala 9:92]
  reg [31:0] _RAND_631;
  reg [7:0] in_rt_wt_data_d_1_116; // @[retiming.scala 9:92]
  reg [31:0] _RAND_632;
  reg [7:0] in_rt_wt_data_d_1_117; // @[retiming.scala 9:92]
  reg [31:0] _RAND_633;
  reg [7:0] in_rt_wt_data_d_1_118; // @[retiming.scala 9:92]
  reg [31:0] _RAND_634;
  reg [7:0] in_rt_wt_data_d_1_119; // @[retiming.scala 9:92]
  reg [31:0] _RAND_635;
  reg [7:0] in_rt_wt_data_d_1_120; // @[retiming.scala 9:92]
  reg [31:0] _RAND_636;
  reg [7:0] in_rt_wt_data_d_1_121; // @[retiming.scala 9:92]
  reg [31:0] _RAND_637;
  reg [7:0] in_rt_wt_data_d_1_122; // @[retiming.scala 9:92]
  reg [31:0] _RAND_638;
  reg [7:0] in_rt_wt_data_d_1_123; // @[retiming.scala 9:92]
  reg [31:0] _RAND_639;
  reg [7:0] in_rt_wt_data_d_1_124; // @[retiming.scala 9:92]
  reg [31:0] _RAND_640;
  reg [7:0] in_rt_wt_data_d_1_125; // @[retiming.scala 9:92]
  reg [31:0] _RAND_641;
  reg [7:0] in_rt_wt_data_d_1_126; // @[retiming.scala 9:92]
  reg [31:0] _RAND_642;
  reg [7:0] in_rt_wt_data_d_1_127; // @[retiming.scala 9:92]
  reg [31:0] _RAND_643;
  reg [7:0] in_rt_wt_data_d_2_0; // @[retiming.scala 9:92]
  reg [31:0] _RAND_644;
  reg [7:0] in_rt_wt_data_d_2_1; // @[retiming.scala 9:92]
  reg [31:0] _RAND_645;
  reg [7:0] in_rt_wt_data_d_2_2; // @[retiming.scala 9:92]
  reg [31:0] _RAND_646;
  reg [7:0] in_rt_wt_data_d_2_3; // @[retiming.scala 9:92]
  reg [31:0] _RAND_647;
  reg [7:0] in_rt_wt_data_d_2_4; // @[retiming.scala 9:92]
  reg [31:0] _RAND_648;
  reg [7:0] in_rt_wt_data_d_2_5; // @[retiming.scala 9:92]
  reg [31:0] _RAND_649;
  reg [7:0] in_rt_wt_data_d_2_6; // @[retiming.scala 9:92]
  reg [31:0] _RAND_650;
  reg [7:0] in_rt_wt_data_d_2_7; // @[retiming.scala 9:92]
  reg [31:0] _RAND_651;
  reg [7:0] in_rt_wt_data_d_2_8; // @[retiming.scala 9:92]
  reg [31:0] _RAND_652;
  reg [7:0] in_rt_wt_data_d_2_9; // @[retiming.scala 9:92]
  reg [31:0] _RAND_653;
  reg [7:0] in_rt_wt_data_d_2_10; // @[retiming.scala 9:92]
  reg [31:0] _RAND_654;
  reg [7:0] in_rt_wt_data_d_2_11; // @[retiming.scala 9:92]
  reg [31:0] _RAND_655;
  reg [7:0] in_rt_wt_data_d_2_12; // @[retiming.scala 9:92]
  reg [31:0] _RAND_656;
  reg [7:0] in_rt_wt_data_d_2_13; // @[retiming.scala 9:92]
  reg [31:0] _RAND_657;
  reg [7:0] in_rt_wt_data_d_2_14; // @[retiming.scala 9:92]
  reg [31:0] _RAND_658;
  reg [7:0] in_rt_wt_data_d_2_15; // @[retiming.scala 9:92]
  reg [31:0] _RAND_659;
  reg [7:0] in_rt_wt_data_d_2_16; // @[retiming.scala 9:92]
  reg [31:0] _RAND_660;
  reg [7:0] in_rt_wt_data_d_2_17; // @[retiming.scala 9:92]
  reg [31:0] _RAND_661;
  reg [7:0] in_rt_wt_data_d_2_18; // @[retiming.scala 9:92]
  reg [31:0] _RAND_662;
  reg [7:0] in_rt_wt_data_d_2_19; // @[retiming.scala 9:92]
  reg [31:0] _RAND_663;
  reg [7:0] in_rt_wt_data_d_2_20; // @[retiming.scala 9:92]
  reg [31:0] _RAND_664;
  reg [7:0] in_rt_wt_data_d_2_21; // @[retiming.scala 9:92]
  reg [31:0] _RAND_665;
  reg [7:0] in_rt_wt_data_d_2_22; // @[retiming.scala 9:92]
  reg [31:0] _RAND_666;
  reg [7:0] in_rt_wt_data_d_2_23; // @[retiming.scala 9:92]
  reg [31:0] _RAND_667;
  reg [7:0] in_rt_wt_data_d_2_24; // @[retiming.scala 9:92]
  reg [31:0] _RAND_668;
  reg [7:0] in_rt_wt_data_d_2_25; // @[retiming.scala 9:92]
  reg [31:0] _RAND_669;
  reg [7:0] in_rt_wt_data_d_2_26; // @[retiming.scala 9:92]
  reg [31:0] _RAND_670;
  reg [7:0] in_rt_wt_data_d_2_27; // @[retiming.scala 9:92]
  reg [31:0] _RAND_671;
  reg [7:0] in_rt_wt_data_d_2_28; // @[retiming.scala 9:92]
  reg [31:0] _RAND_672;
  reg [7:0] in_rt_wt_data_d_2_29; // @[retiming.scala 9:92]
  reg [31:0] _RAND_673;
  reg [7:0] in_rt_wt_data_d_2_30; // @[retiming.scala 9:92]
  reg [31:0] _RAND_674;
  reg [7:0] in_rt_wt_data_d_2_31; // @[retiming.scala 9:92]
  reg [31:0] _RAND_675;
  reg [7:0] in_rt_wt_data_d_2_32; // @[retiming.scala 9:92]
  reg [31:0] _RAND_676;
  reg [7:0] in_rt_wt_data_d_2_33; // @[retiming.scala 9:92]
  reg [31:0] _RAND_677;
  reg [7:0] in_rt_wt_data_d_2_34; // @[retiming.scala 9:92]
  reg [31:0] _RAND_678;
  reg [7:0] in_rt_wt_data_d_2_35; // @[retiming.scala 9:92]
  reg [31:0] _RAND_679;
  reg [7:0] in_rt_wt_data_d_2_36; // @[retiming.scala 9:92]
  reg [31:0] _RAND_680;
  reg [7:0] in_rt_wt_data_d_2_37; // @[retiming.scala 9:92]
  reg [31:0] _RAND_681;
  reg [7:0] in_rt_wt_data_d_2_38; // @[retiming.scala 9:92]
  reg [31:0] _RAND_682;
  reg [7:0] in_rt_wt_data_d_2_39; // @[retiming.scala 9:92]
  reg [31:0] _RAND_683;
  reg [7:0] in_rt_wt_data_d_2_40; // @[retiming.scala 9:92]
  reg [31:0] _RAND_684;
  reg [7:0] in_rt_wt_data_d_2_41; // @[retiming.scala 9:92]
  reg [31:0] _RAND_685;
  reg [7:0] in_rt_wt_data_d_2_42; // @[retiming.scala 9:92]
  reg [31:0] _RAND_686;
  reg [7:0] in_rt_wt_data_d_2_43; // @[retiming.scala 9:92]
  reg [31:0] _RAND_687;
  reg [7:0] in_rt_wt_data_d_2_44; // @[retiming.scala 9:92]
  reg [31:0] _RAND_688;
  reg [7:0] in_rt_wt_data_d_2_45; // @[retiming.scala 9:92]
  reg [31:0] _RAND_689;
  reg [7:0] in_rt_wt_data_d_2_46; // @[retiming.scala 9:92]
  reg [31:0] _RAND_690;
  reg [7:0] in_rt_wt_data_d_2_47; // @[retiming.scala 9:92]
  reg [31:0] _RAND_691;
  reg [7:0] in_rt_wt_data_d_2_48; // @[retiming.scala 9:92]
  reg [31:0] _RAND_692;
  reg [7:0] in_rt_wt_data_d_2_49; // @[retiming.scala 9:92]
  reg [31:0] _RAND_693;
  reg [7:0] in_rt_wt_data_d_2_50; // @[retiming.scala 9:92]
  reg [31:0] _RAND_694;
  reg [7:0] in_rt_wt_data_d_2_51; // @[retiming.scala 9:92]
  reg [31:0] _RAND_695;
  reg [7:0] in_rt_wt_data_d_2_52; // @[retiming.scala 9:92]
  reg [31:0] _RAND_696;
  reg [7:0] in_rt_wt_data_d_2_53; // @[retiming.scala 9:92]
  reg [31:0] _RAND_697;
  reg [7:0] in_rt_wt_data_d_2_54; // @[retiming.scala 9:92]
  reg [31:0] _RAND_698;
  reg [7:0] in_rt_wt_data_d_2_55; // @[retiming.scala 9:92]
  reg [31:0] _RAND_699;
  reg [7:0] in_rt_wt_data_d_2_56; // @[retiming.scala 9:92]
  reg [31:0] _RAND_700;
  reg [7:0] in_rt_wt_data_d_2_57; // @[retiming.scala 9:92]
  reg [31:0] _RAND_701;
  reg [7:0] in_rt_wt_data_d_2_58; // @[retiming.scala 9:92]
  reg [31:0] _RAND_702;
  reg [7:0] in_rt_wt_data_d_2_59; // @[retiming.scala 9:92]
  reg [31:0] _RAND_703;
  reg [7:0] in_rt_wt_data_d_2_60; // @[retiming.scala 9:92]
  reg [31:0] _RAND_704;
  reg [7:0] in_rt_wt_data_d_2_61; // @[retiming.scala 9:92]
  reg [31:0] _RAND_705;
  reg [7:0] in_rt_wt_data_d_2_62; // @[retiming.scala 9:92]
  reg [31:0] _RAND_706;
  reg [7:0] in_rt_wt_data_d_2_63; // @[retiming.scala 9:92]
  reg [31:0] _RAND_707;
  reg [7:0] in_rt_wt_data_d_2_64; // @[retiming.scala 9:92]
  reg [31:0] _RAND_708;
  reg [7:0] in_rt_wt_data_d_2_65; // @[retiming.scala 9:92]
  reg [31:0] _RAND_709;
  reg [7:0] in_rt_wt_data_d_2_66; // @[retiming.scala 9:92]
  reg [31:0] _RAND_710;
  reg [7:0] in_rt_wt_data_d_2_67; // @[retiming.scala 9:92]
  reg [31:0] _RAND_711;
  reg [7:0] in_rt_wt_data_d_2_68; // @[retiming.scala 9:92]
  reg [31:0] _RAND_712;
  reg [7:0] in_rt_wt_data_d_2_69; // @[retiming.scala 9:92]
  reg [31:0] _RAND_713;
  reg [7:0] in_rt_wt_data_d_2_70; // @[retiming.scala 9:92]
  reg [31:0] _RAND_714;
  reg [7:0] in_rt_wt_data_d_2_71; // @[retiming.scala 9:92]
  reg [31:0] _RAND_715;
  reg [7:0] in_rt_wt_data_d_2_72; // @[retiming.scala 9:92]
  reg [31:0] _RAND_716;
  reg [7:0] in_rt_wt_data_d_2_73; // @[retiming.scala 9:92]
  reg [31:0] _RAND_717;
  reg [7:0] in_rt_wt_data_d_2_74; // @[retiming.scala 9:92]
  reg [31:0] _RAND_718;
  reg [7:0] in_rt_wt_data_d_2_75; // @[retiming.scala 9:92]
  reg [31:0] _RAND_719;
  reg [7:0] in_rt_wt_data_d_2_76; // @[retiming.scala 9:92]
  reg [31:0] _RAND_720;
  reg [7:0] in_rt_wt_data_d_2_77; // @[retiming.scala 9:92]
  reg [31:0] _RAND_721;
  reg [7:0] in_rt_wt_data_d_2_78; // @[retiming.scala 9:92]
  reg [31:0] _RAND_722;
  reg [7:0] in_rt_wt_data_d_2_79; // @[retiming.scala 9:92]
  reg [31:0] _RAND_723;
  reg [7:0] in_rt_wt_data_d_2_80; // @[retiming.scala 9:92]
  reg [31:0] _RAND_724;
  reg [7:0] in_rt_wt_data_d_2_81; // @[retiming.scala 9:92]
  reg [31:0] _RAND_725;
  reg [7:0] in_rt_wt_data_d_2_82; // @[retiming.scala 9:92]
  reg [31:0] _RAND_726;
  reg [7:0] in_rt_wt_data_d_2_83; // @[retiming.scala 9:92]
  reg [31:0] _RAND_727;
  reg [7:0] in_rt_wt_data_d_2_84; // @[retiming.scala 9:92]
  reg [31:0] _RAND_728;
  reg [7:0] in_rt_wt_data_d_2_85; // @[retiming.scala 9:92]
  reg [31:0] _RAND_729;
  reg [7:0] in_rt_wt_data_d_2_86; // @[retiming.scala 9:92]
  reg [31:0] _RAND_730;
  reg [7:0] in_rt_wt_data_d_2_87; // @[retiming.scala 9:92]
  reg [31:0] _RAND_731;
  reg [7:0] in_rt_wt_data_d_2_88; // @[retiming.scala 9:92]
  reg [31:0] _RAND_732;
  reg [7:0] in_rt_wt_data_d_2_89; // @[retiming.scala 9:92]
  reg [31:0] _RAND_733;
  reg [7:0] in_rt_wt_data_d_2_90; // @[retiming.scala 9:92]
  reg [31:0] _RAND_734;
  reg [7:0] in_rt_wt_data_d_2_91; // @[retiming.scala 9:92]
  reg [31:0] _RAND_735;
  reg [7:0] in_rt_wt_data_d_2_92; // @[retiming.scala 9:92]
  reg [31:0] _RAND_736;
  reg [7:0] in_rt_wt_data_d_2_93; // @[retiming.scala 9:92]
  reg [31:0] _RAND_737;
  reg [7:0] in_rt_wt_data_d_2_94; // @[retiming.scala 9:92]
  reg [31:0] _RAND_738;
  reg [7:0] in_rt_wt_data_d_2_95; // @[retiming.scala 9:92]
  reg [31:0] _RAND_739;
  reg [7:0] in_rt_wt_data_d_2_96; // @[retiming.scala 9:92]
  reg [31:0] _RAND_740;
  reg [7:0] in_rt_wt_data_d_2_97; // @[retiming.scala 9:92]
  reg [31:0] _RAND_741;
  reg [7:0] in_rt_wt_data_d_2_98; // @[retiming.scala 9:92]
  reg [31:0] _RAND_742;
  reg [7:0] in_rt_wt_data_d_2_99; // @[retiming.scala 9:92]
  reg [31:0] _RAND_743;
  reg [7:0] in_rt_wt_data_d_2_100; // @[retiming.scala 9:92]
  reg [31:0] _RAND_744;
  reg [7:0] in_rt_wt_data_d_2_101; // @[retiming.scala 9:92]
  reg [31:0] _RAND_745;
  reg [7:0] in_rt_wt_data_d_2_102; // @[retiming.scala 9:92]
  reg [31:0] _RAND_746;
  reg [7:0] in_rt_wt_data_d_2_103; // @[retiming.scala 9:92]
  reg [31:0] _RAND_747;
  reg [7:0] in_rt_wt_data_d_2_104; // @[retiming.scala 9:92]
  reg [31:0] _RAND_748;
  reg [7:0] in_rt_wt_data_d_2_105; // @[retiming.scala 9:92]
  reg [31:0] _RAND_749;
  reg [7:0] in_rt_wt_data_d_2_106; // @[retiming.scala 9:92]
  reg [31:0] _RAND_750;
  reg [7:0] in_rt_wt_data_d_2_107; // @[retiming.scala 9:92]
  reg [31:0] _RAND_751;
  reg [7:0] in_rt_wt_data_d_2_108; // @[retiming.scala 9:92]
  reg [31:0] _RAND_752;
  reg [7:0] in_rt_wt_data_d_2_109; // @[retiming.scala 9:92]
  reg [31:0] _RAND_753;
  reg [7:0] in_rt_wt_data_d_2_110; // @[retiming.scala 9:92]
  reg [31:0] _RAND_754;
  reg [7:0] in_rt_wt_data_d_2_111; // @[retiming.scala 9:92]
  reg [31:0] _RAND_755;
  reg [7:0] in_rt_wt_data_d_2_112; // @[retiming.scala 9:92]
  reg [31:0] _RAND_756;
  reg [7:0] in_rt_wt_data_d_2_113; // @[retiming.scala 9:92]
  reg [31:0] _RAND_757;
  reg [7:0] in_rt_wt_data_d_2_114; // @[retiming.scala 9:92]
  reg [31:0] _RAND_758;
  reg [7:0] in_rt_wt_data_d_2_115; // @[retiming.scala 9:92]
  reg [31:0] _RAND_759;
  reg [7:0] in_rt_wt_data_d_2_116; // @[retiming.scala 9:92]
  reg [31:0] _RAND_760;
  reg [7:0] in_rt_wt_data_d_2_117; // @[retiming.scala 9:92]
  reg [31:0] _RAND_761;
  reg [7:0] in_rt_wt_data_d_2_118; // @[retiming.scala 9:92]
  reg [31:0] _RAND_762;
  reg [7:0] in_rt_wt_data_d_2_119; // @[retiming.scala 9:92]
  reg [31:0] _RAND_763;
  reg [7:0] in_rt_wt_data_d_2_120; // @[retiming.scala 9:92]
  reg [31:0] _RAND_764;
  reg [7:0] in_rt_wt_data_d_2_121; // @[retiming.scala 9:92]
  reg [31:0] _RAND_765;
  reg [7:0] in_rt_wt_data_d_2_122; // @[retiming.scala 9:92]
  reg [31:0] _RAND_766;
  reg [7:0] in_rt_wt_data_d_2_123; // @[retiming.scala 9:92]
  reg [31:0] _RAND_767;
  reg [7:0] in_rt_wt_data_d_2_124; // @[retiming.scala 9:92]
  reg [31:0] _RAND_768;
  reg [7:0] in_rt_wt_data_d_2_125; // @[retiming.scala 9:92]
  reg [31:0] _RAND_769;
  reg [7:0] in_rt_wt_data_d_2_126; // @[retiming.scala 9:92]
  reg [31:0] _RAND_770;
  reg [7:0] in_rt_wt_data_d_2_127; // @[retiming.scala 9:92]
  reg [31:0] _RAND_771;
  reg  in_rt_wt_mask_d_1_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_772;
  reg  in_rt_wt_mask_d_1_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_773;
  reg  in_rt_wt_mask_d_1_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_774;
  reg  in_rt_wt_mask_d_1_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_775;
  reg  in_rt_wt_mask_d_1_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_776;
  reg  in_rt_wt_mask_d_1_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_777;
  reg  in_rt_wt_mask_d_1_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_778;
  reg  in_rt_wt_mask_d_1_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_779;
  reg  in_rt_wt_mask_d_1_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_780;
  reg  in_rt_wt_mask_d_1_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_781;
  reg  in_rt_wt_mask_d_1_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_782;
  reg  in_rt_wt_mask_d_1_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_783;
  reg  in_rt_wt_mask_d_1_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_784;
  reg  in_rt_wt_mask_d_1_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_785;
  reg  in_rt_wt_mask_d_1_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_786;
  reg  in_rt_wt_mask_d_1_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_787;
  reg  in_rt_wt_mask_d_1_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_788;
  reg  in_rt_wt_mask_d_1_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_789;
  reg  in_rt_wt_mask_d_1_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_790;
  reg  in_rt_wt_mask_d_1_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_791;
  reg  in_rt_wt_mask_d_1_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_792;
  reg  in_rt_wt_mask_d_1_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_793;
  reg  in_rt_wt_mask_d_1_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_794;
  reg  in_rt_wt_mask_d_1_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_795;
  reg  in_rt_wt_mask_d_1_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_796;
  reg  in_rt_wt_mask_d_1_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_797;
  reg  in_rt_wt_mask_d_1_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_798;
  reg  in_rt_wt_mask_d_1_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_799;
  reg  in_rt_wt_mask_d_1_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_800;
  reg  in_rt_wt_mask_d_1_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_801;
  reg  in_rt_wt_mask_d_1_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_802;
  reg  in_rt_wt_mask_d_1_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_803;
  reg  in_rt_wt_mask_d_1_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_804;
  reg  in_rt_wt_mask_d_1_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_805;
  reg  in_rt_wt_mask_d_1_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_806;
  reg  in_rt_wt_mask_d_1_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_807;
  reg  in_rt_wt_mask_d_1_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_808;
  reg  in_rt_wt_mask_d_1_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_809;
  reg  in_rt_wt_mask_d_1_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_810;
  reg  in_rt_wt_mask_d_1_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_811;
  reg  in_rt_wt_mask_d_1_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_812;
  reg  in_rt_wt_mask_d_1_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_813;
  reg  in_rt_wt_mask_d_1_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_814;
  reg  in_rt_wt_mask_d_1_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_815;
  reg  in_rt_wt_mask_d_1_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_816;
  reg  in_rt_wt_mask_d_1_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_817;
  reg  in_rt_wt_mask_d_1_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_818;
  reg  in_rt_wt_mask_d_1_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_819;
  reg  in_rt_wt_mask_d_1_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_820;
  reg  in_rt_wt_mask_d_1_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_821;
  reg  in_rt_wt_mask_d_1_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_822;
  reg  in_rt_wt_mask_d_1_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_823;
  reg  in_rt_wt_mask_d_1_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_824;
  reg  in_rt_wt_mask_d_1_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_825;
  reg  in_rt_wt_mask_d_1_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_826;
  reg  in_rt_wt_mask_d_1_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_827;
  reg  in_rt_wt_mask_d_1_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_828;
  reg  in_rt_wt_mask_d_1_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_829;
  reg  in_rt_wt_mask_d_1_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_830;
  reg  in_rt_wt_mask_d_1_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_831;
  reg  in_rt_wt_mask_d_1_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_832;
  reg  in_rt_wt_mask_d_1_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_833;
  reg  in_rt_wt_mask_d_1_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_834;
  reg  in_rt_wt_mask_d_1_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_835;
  reg  in_rt_wt_mask_d_1_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_836;
  reg  in_rt_wt_mask_d_1_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_837;
  reg  in_rt_wt_mask_d_1_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_838;
  reg  in_rt_wt_mask_d_1_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_839;
  reg  in_rt_wt_mask_d_1_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_840;
  reg  in_rt_wt_mask_d_1_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_841;
  reg  in_rt_wt_mask_d_1_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_842;
  reg  in_rt_wt_mask_d_1_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_843;
  reg  in_rt_wt_mask_d_1_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_844;
  reg  in_rt_wt_mask_d_1_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_845;
  reg  in_rt_wt_mask_d_1_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_846;
  reg  in_rt_wt_mask_d_1_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_847;
  reg  in_rt_wt_mask_d_1_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_848;
  reg  in_rt_wt_mask_d_1_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_849;
  reg  in_rt_wt_mask_d_1_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_850;
  reg  in_rt_wt_mask_d_1_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_851;
  reg  in_rt_wt_mask_d_1_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_852;
  reg  in_rt_wt_mask_d_1_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_853;
  reg  in_rt_wt_mask_d_1_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_854;
  reg  in_rt_wt_mask_d_1_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_855;
  reg  in_rt_wt_mask_d_1_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_856;
  reg  in_rt_wt_mask_d_1_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_857;
  reg  in_rt_wt_mask_d_1_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_858;
  reg  in_rt_wt_mask_d_1_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_859;
  reg  in_rt_wt_mask_d_1_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_860;
  reg  in_rt_wt_mask_d_1_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_861;
  reg  in_rt_wt_mask_d_1_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_862;
  reg  in_rt_wt_mask_d_1_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_863;
  reg  in_rt_wt_mask_d_1_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_864;
  reg  in_rt_wt_mask_d_1_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_865;
  reg  in_rt_wt_mask_d_1_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_866;
  reg  in_rt_wt_mask_d_1_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_867;
  reg  in_rt_wt_mask_d_1_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_868;
  reg  in_rt_wt_mask_d_1_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_869;
  reg  in_rt_wt_mask_d_1_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_870;
  reg  in_rt_wt_mask_d_1_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_871;
  reg  in_rt_wt_mask_d_1_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_872;
  reg  in_rt_wt_mask_d_1_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_873;
  reg  in_rt_wt_mask_d_1_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_874;
  reg  in_rt_wt_mask_d_1_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_875;
  reg  in_rt_wt_mask_d_1_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_876;
  reg  in_rt_wt_mask_d_1_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_877;
  reg  in_rt_wt_mask_d_1_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_878;
  reg  in_rt_wt_mask_d_1_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_879;
  reg  in_rt_wt_mask_d_1_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_880;
  reg  in_rt_wt_mask_d_1_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_881;
  reg  in_rt_wt_mask_d_1_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_882;
  reg  in_rt_wt_mask_d_1_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_883;
  reg  in_rt_wt_mask_d_1_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_884;
  reg  in_rt_wt_mask_d_1_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_885;
  reg  in_rt_wt_mask_d_1_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_886;
  reg  in_rt_wt_mask_d_1_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_887;
  reg  in_rt_wt_mask_d_1_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_888;
  reg  in_rt_wt_mask_d_1_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_889;
  reg  in_rt_wt_mask_d_1_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_890;
  reg  in_rt_wt_mask_d_1_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_891;
  reg  in_rt_wt_mask_d_1_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_892;
  reg  in_rt_wt_mask_d_1_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_893;
  reg  in_rt_wt_mask_d_1_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_894;
  reg  in_rt_wt_mask_d_1_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_895;
  reg  in_rt_wt_mask_d_1_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_896;
  reg  in_rt_wt_mask_d_1_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_897;
  reg  in_rt_wt_mask_d_1_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_898;
  reg  in_rt_wt_mask_d_1_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_899;
  reg  in_rt_wt_mask_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_900;
  reg  in_rt_wt_mask_d_2_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_901;
  reg  in_rt_wt_mask_d_2_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_902;
  reg  in_rt_wt_mask_d_2_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_903;
  reg  in_rt_wt_mask_d_2_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_904;
  reg  in_rt_wt_mask_d_2_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_905;
  reg  in_rt_wt_mask_d_2_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_906;
  reg  in_rt_wt_mask_d_2_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_907;
  reg  in_rt_wt_mask_d_2_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_908;
  reg  in_rt_wt_mask_d_2_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_909;
  reg  in_rt_wt_mask_d_2_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_910;
  reg  in_rt_wt_mask_d_2_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_911;
  reg  in_rt_wt_mask_d_2_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_912;
  reg  in_rt_wt_mask_d_2_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_913;
  reg  in_rt_wt_mask_d_2_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_914;
  reg  in_rt_wt_mask_d_2_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_915;
  reg  in_rt_wt_mask_d_2_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_916;
  reg  in_rt_wt_mask_d_2_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_917;
  reg  in_rt_wt_mask_d_2_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_918;
  reg  in_rt_wt_mask_d_2_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_919;
  reg  in_rt_wt_mask_d_2_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_920;
  reg  in_rt_wt_mask_d_2_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_921;
  reg  in_rt_wt_mask_d_2_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_922;
  reg  in_rt_wt_mask_d_2_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_923;
  reg  in_rt_wt_mask_d_2_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_924;
  reg  in_rt_wt_mask_d_2_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_925;
  reg  in_rt_wt_mask_d_2_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_926;
  reg  in_rt_wt_mask_d_2_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_927;
  reg  in_rt_wt_mask_d_2_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_928;
  reg  in_rt_wt_mask_d_2_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_929;
  reg  in_rt_wt_mask_d_2_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_930;
  reg  in_rt_wt_mask_d_2_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_931;
  reg  in_rt_wt_mask_d_2_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_932;
  reg  in_rt_wt_mask_d_2_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_933;
  reg  in_rt_wt_mask_d_2_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_934;
  reg  in_rt_wt_mask_d_2_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_935;
  reg  in_rt_wt_mask_d_2_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_936;
  reg  in_rt_wt_mask_d_2_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_937;
  reg  in_rt_wt_mask_d_2_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_938;
  reg  in_rt_wt_mask_d_2_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_939;
  reg  in_rt_wt_mask_d_2_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_940;
  reg  in_rt_wt_mask_d_2_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_941;
  reg  in_rt_wt_mask_d_2_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_942;
  reg  in_rt_wt_mask_d_2_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_943;
  reg  in_rt_wt_mask_d_2_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_944;
  reg  in_rt_wt_mask_d_2_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_945;
  reg  in_rt_wt_mask_d_2_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_946;
  reg  in_rt_wt_mask_d_2_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_947;
  reg  in_rt_wt_mask_d_2_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_948;
  reg  in_rt_wt_mask_d_2_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_949;
  reg  in_rt_wt_mask_d_2_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_950;
  reg  in_rt_wt_mask_d_2_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_951;
  reg  in_rt_wt_mask_d_2_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_952;
  reg  in_rt_wt_mask_d_2_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_953;
  reg  in_rt_wt_mask_d_2_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_954;
  reg  in_rt_wt_mask_d_2_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_955;
  reg  in_rt_wt_mask_d_2_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_956;
  reg  in_rt_wt_mask_d_2_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_957;
  reg  in_rt_wt_mask_d_2_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_958;
  reg  in_rt_wt_mask_d_2_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_959;
  reg  in_rt_wt_mask_d_2_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_960;
  reg  in_rt_wt_mask_d_2_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_961;
  reg  in_rt_wt_mask_d_2_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_962;
  reg  in_rt_wt_mask_d_2_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_963;
  reg  in_rt_wt_mask_d_2_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_964;
  reg  in_rt_wt_mask_d_2_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_965;
  reg  in_rt_wt_mask_d_2_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_966;
  reg  in_rt_wt_mask_d_2_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_967;
  reg  in_rt_wt_mask_d_2_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_968;
  reg  in_rt_wt_mask_d_2_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_969;
  reg  in_rt_wt_mask_d_2_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_970;
  reg  in_rt_wt_mask_d_2_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_971;
  reg  in_rt_wt_mask_d_2_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_972;
  reg  in_rt_wt_mask_d_2_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_973;
  reg  in_rt_wt_mask_d_2_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_974;
  reg  in_rt_wt_mask_d_2_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_975;
  reg  in_rt_wt_mask_d_2_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_976;
  reg  in_rt_wt_mask_d_2_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_977;
  reg  in_rt_wt_mask_d_2_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_978;
  reg  in_rt_wt_mask_d_2_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_979;
  reg  in_rt_wt_mask_d_2_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_980;
  reg  in_rt_wt_mask_d_2_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_981;
  reg  in_rt_wt_mask_d_2_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_982;
  reg  in_rt_wt_mask_d_2_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_983;
  reg  in_rt_wt_mask_d_2_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_984;
  reg  in_rt_wt_mask_d_2_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_985;
  reg  in_rt_wt_mask_d_2_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_986;
  reg  in_rt_wt_mask_d_2_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_987;
  reg  in_rt_wt_mask_d_2_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_988;
  reg  in_rt_wt_mask_d_2_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_989;
  reg  in_rt_wt_mask_d_2_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_990;
  reg  in_rt_wt_mask_d_2_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_991;
  reg  in_rt_wt_mask_d_2_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_992;
  reg  in_rt_wt_mask_d_2_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_993;
  reg  in_rt_wt_mask_d_2_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_994;
  reg  in_rt_wt_mask_d_2_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_995;
  reg  in_rt_wt_mask_d_2_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_996;
  reg  in_rt_wt_mask_d_2_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_997;
  reg  in_rt_wt_mask_d_2_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_998;
  reg  in_rt_wt_mask_d_2_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_999;
  reg  in_rt_wt_mask_d_2_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1000;
  reg  in_rt_wt_mask_d_2_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1001;
  reg  in_rt_wt_mask_d_2_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1002;
  reg  in_rt_wt_mask_d_2_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1003;
  reg  in_rt_wt_mask_d_2_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1004;
  reg  in_rt_wt_mask_d_2_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1005;
  reg  in_rt_wt_mask_d_2_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1006;
  reg  in_rt_wt_mask_d_2_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1007;
  reg  in_rt_wt_mask_d_2_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1008;
  reg  in_rt_wt_mask_d_2_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1009;
  reg  in_rt_wt_mask_d_2_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1010;
  reg  in_rt_wt_mask_d_2_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1011;
  reg  in_rt_wt_mask_d_2_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1012;
  reg  in_rt_wt_mask_d_2_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1013;
  reg  in_rt_wt_mask_d_2_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1014;
  reg  in_rt_wt_mask_d_2_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1015;
  reg  in_rt_wt_mask_d_2_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1016;
  reg  in_rt_wt_mask_d_2_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1017;
  reg  in_rt_wt_mask_d_2_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1018;
  reg  in_rt_wt_mask_d_2_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1019;
  reg  in_rt_wt_mask_d_2_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1020;
  reg  in_rt_wt_mask_d_2_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1021;
  reg  in_rt_wt_mask_d_2_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1022;
  reg  in_rt_wt_mask_d_2_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1023;
  reg  in_rt_wt_mask_d_2_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1024;
  reg  in_rt_wt_mask_d_2_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1025;
  reg  in_rt_wt_mask_d_2_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1026;
  reg  in_rt_wt_mask_d_2_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 69:70]
  reg [31:0] _RAND_1027;
  reg  in_rt_wt_pvld_d_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 71:70]
  reg [31:0] _RAND_1028;
  reg  in_rt_wt_pvld_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 71:70]
  reg [31:0] _RAND_1029;
  reg  in_rt_wt_sel_d_1_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 73:70]
  reg [31:0] _RAND_1030;
  reg  in_rt_wt_sel_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 73:70]
  reg [31:0] _RAND_1031;
  wire  _T_6928; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:33]
  wire  _GEN_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire [8:0] _GEN_128; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _T_6929; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:32]
  wire  _GEN_129; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_130; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_131; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_132; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_133; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_134; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_135; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_136; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_137; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_138; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_139; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_140; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_141; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_142; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_143; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_144; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_145; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_146; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_147; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_148; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_149; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_150; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_151; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_152; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_153; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_154; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_155; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_156; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_157; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_158; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_159; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_160; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_161; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_162; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_163; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_164; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_165; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_166; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_167; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_168; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_169; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_170; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_171; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_172; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_173; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_174; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_175; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_176; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_177; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_178; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_179; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_180; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_181; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_182; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_183; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_184; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_185; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_186; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_187; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_188; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_189; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_190; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_191; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_192; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_193; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_194; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_195; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_196; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_197; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_198; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_199; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_200; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_201; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_202; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_203; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_204; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_205; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_206; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_207; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_208; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_209; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_210; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_211; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_212; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_213; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_214; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_215; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_216; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_217; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_218; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_219; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_220; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_221; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_222; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_223; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_224; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_225; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_226; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_227; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_228; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_229; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_230; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_231; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_232; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_233; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_234; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_235; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_236; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_237; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_238; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_239; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_240; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_241; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_242; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_243; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_244; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_245; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_246; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_247; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_248; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_249; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_250; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_251; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_252; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_253; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_254; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_255; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_256; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_257; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _T_6930; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:33]
  wire  _GEN_514; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_515; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_516; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_517; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_518; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_519; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_520; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_521; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_522; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_523; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_524; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_525; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_526; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_527; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_528; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_529; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_530; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_531; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_532; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_533; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_534; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_535; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_536; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_537; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_538; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_539; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_540; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_541; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_542; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_543; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_544; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_545; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_546; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_547; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_548; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_549; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_550; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_551; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_552; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_553; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_554; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_555; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_556; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_557; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_558; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_559; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_560; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_561; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_562; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_563; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_564; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_565; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_566; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_567; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_568; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_569; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_570; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_571; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_572; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_573; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_574; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_575; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_576; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_577; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_578; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_579; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_580; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_581; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_582; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_583; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_584; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_585; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_586; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_587; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_588; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_589; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_590; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_591; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_592; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_593; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_594; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_595; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_596; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_597; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_598; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_599; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_600; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_601; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_602; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_603; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_604; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_605; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_606; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_607; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_608; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_609; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_610; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_611; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_612; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_613; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_614; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_615; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_616; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_617; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_618; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_619; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_620; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_621; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_622; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_623; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_624; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_625; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_626; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_627; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_628; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_629; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_630; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_631; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_632; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_633; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_634; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_635; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_636; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_637; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_638; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_639; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_640; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _GEN_641; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire [8:0] _GEN_642; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  wire  _T_6931; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:32]
  wire  _GEN_643; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_644; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_645; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_646; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_647; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_648; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_649; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_650; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_651; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_652; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_653; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_654; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_655; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_656; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_657; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_658; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_659; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_660; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_661; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_662; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_663; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_664; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_665; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_666; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_667; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_668; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_669; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_670; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_671; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_672; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_673; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_674; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_675; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_676; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_677; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_678; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_679; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_680; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_681; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_682; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_683; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_684; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_685; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_686; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_687; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_688; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_689; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_690; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_691; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_692; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_693; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_694; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_695; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_696; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_697; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_698; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_699; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_700; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_701; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_702; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_703; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_704; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_705; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_706; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_707; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_708; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_709; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_710; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_711; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_712; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_713; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_714; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_715; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_716; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_717; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_718; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_719; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_720; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_721; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_722; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_723; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_724; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_725; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_726; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_727; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_728; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_729; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_730; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_731; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_732; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_733; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_734; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_735; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_736; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_737; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_738; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_739; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_740; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_741; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_742; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_743; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_744; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_745; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_746; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_747; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_748; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_749; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_750; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_751; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_752; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_753; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_754; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_755; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_756; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_757; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_758; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_759; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_760; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_761; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_762; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_763; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_764; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_765; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_766; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_767; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_768; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_769; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_770; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  wire  _GEN_771; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _T_6928 = io_sc2mac_dat_pvld | in_rt_dat_pvld_d_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:33]
  assign _GEN_0 = _T_6928 ? io_sc2mac_dat_mask_0 : in_rt_dat_mask_d_1_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_1 = _T_6928 ? io_sc2mac_dat_mask_1 : in_rt_dat_mask_d_1_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_2 = _T_6928 ? io_sc2mac_dat_mask_2 : in_rt_dat_mask_d_1_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_3 = _T_6928 ? io_sc2mac_dat_mask_3 : in_rt_dat_mask_d_1_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_4 = _T_6928 ? io_sc2mac_dat_mask_4 : in_rt_dat_mask_d_1_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_5 = _T_6928 ? io_sc2mac_dat_mask_5 : in_rt_dat_mask_d_1_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_6 = _T_6928 ? io_sc2mac_dat_mask_6 : in_rt_dat_mask_d_1_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_7 = _T_6928 ? io_sc2mac_dat_mask_7 : in_rt_dat_mask_d_1_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_8 = _T_6928 ? io_sc2mac_dat_mask_8 : in_rt_dat_mask_d_1_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_9 = _T_6928 ? io_sc2mac_dat_mask_9 : in_rt_dat_mask_d_1_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_10 = _T_6928 ? io_sc2mac_dat_mask_10 : in_rt_dat_mask_d_1_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_11 = _T_6928 ? io_sc2mac_dat_mask_11 : in_rt_dat_mask_d_1_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_12 = _T_6928 ? io_sc2mac_dat_mask_12 : in_rt_dat_mask_d_1_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_13 = _T_6928 ? io_sc2mac_dat_mask_13 : in_rt_dat_mask_d_1_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_14 = _T_6928 ? io_sc2mac_dat_mask_14 : in_rt_dat_mask_d_1_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_15 = _T_6928 ? io_sc2mac_dat_mask_15 : in_rt_dat_mask_d_1_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_16 = _T_6928 ? io_sc2mac_dat_mask_16 : in_rt_dat_mask_d_1_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_17 = _T_6928 ? io_sc2mac_dat_mask_17 : in_rt_dat_mask_d_1_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_18 = _T_6928 ? io_sc2mac_dat_mask_18 : in_rt_dat_mask_d_1_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_19 = _T_6928 ? io_sc2mac_dat_mask_19 : in_rt_dat_mask_d_1_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_20 = _T_6928 ? io_sc2mac_dat_mask_20 : in_rt_dat_mask_d_1_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_21 = _T_6928 ? io_sc2mac_dat_mask_21 : in_rt_dat_mask_d_1_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_22 = _T_6928 ? io_sc2mac_dat_mask_22 : in_rt_dat_mask_d_1_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_23 = _T_6928 ? io_sc2mac_dat_mask_23 : in_rt_dat_mask_d_1_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_24 = _T_6928 ? io_sc2mac_dat_mask_24 : in_rt_dat_mask_d_1_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_25 = _T_6928 ? io_sc2mac_dat_mask_25 : in_rt_dat_mask_d_1_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_26 = _T_6928 ? io_sc2mac_dat_mask_26 : in_rt_dat_mask_d_1_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_27 = _T_6928 ? io_sc2mac_dat_mask_27 : in_rt_dat_mask_d_1_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_28 = _T_6928 ? io_sc2mac_dat_mask_28 : in_rt_dat_mask_d_1_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_29 = _T_6928 ? io_sc2mac_dat_mask_29 : in_rt_dat_mask_d_1_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_30 = _T_6928 ? io_sc2mac_dat_mask_30 : in_rt_dat_mask_d_1_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_31 = _T_6928 ? io_sc2mac_dat_mask_31 : in_rt_dat_mask_d_1_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_32 = _T_6928 ? io_sc2mac_dat_mask_32 : in_rt_dat_mask_d_1_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_33 = _T_6928 ? io_sc2mac_dat_mask_33 : in_rt_dat_mask_d_1_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_34 = _T_6928 ? io_sc2mac_dat_mask_34 : in_rt_dat_mask_d_1_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_35 = _T_6928 ? io_sc2mac_dat_mask_35 : in_rt_dat_mask_d_1_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_36 = _T_6928 ? io_sc2mac_dat_mask_36 : in_rt_dat_mask_d_1_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_37 = _T_6928 ? io_sc2mac_dat_mask_37 : in_rt_dat_mask_d_1_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_38 = _T_6928 ? io_sc2mac_dat_mask_38 : in_rt_dat_mask_d_1_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_39 = _T_6928 ? io_sc2mac_dat_mask_39 : in_rt_dat_mask_d_1_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_40 = _T_6928 ? io_sc2mac_dat_mask_40 : in_rt_dat_mask_d_1_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_41 = _T_6928 ? io_sc2mac_dat_mask_41 : in_rt_dat_mask_d_1_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_42 = _T_6928 ? io_sc2mac_dat_mask_42 : in_rt_dat_mask_d_1_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_43 = _T_6928 ? io_sc2mac_dat_mask_43 : in_rt_dat_mask_d_1_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_44 = _T_6928 ? io_sc2mac_dat_mask_44 : in_rt_dat_mask_d_1_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_45 = _T_6928 ? io_sc2mac_dat_mask_45 : in_rt_dat_mask_d_1_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_46 = _T_6928 ? io_sc2mac_dat_mask_46 : in_rt_dat_mask_d_1_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_47 = _T_6928 ? io_sc2mac_dat_mask_47 : in_rt_dat_mask_d_1_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_48 = _T_6928 ? io_sc2mac_dat_mask_48 : in_rt_dat_mask_d_1_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_49 = _T_6928 ? io_sc2mac_dat_mask_49 : in_rt_dat_mask_d_1_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_50 = _T_6928 ? io_sc2mac_dat_mask_50 : in_rt_dat_mask_d_1_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_51 = _T_6928 ? io_sc2mac_dat_mask_51 : in_rt_dat_mask_d_1_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_52 = _T_6928 ? io_sc2mac_dat_mask_52 : in_rt_dat_mask_d_1_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_53 = _T_6928 ? io_sc2mac_dat_mask_53 : in_rt_dat_mask_d_1_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_54 = _T_6928 ? io_sc2mac_dat_mask_54 : in_rt_dat_mask_d_1_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_55 = _T_6928 ? io_sc2mac_dat_mask_55 : in_rt_dat_mask_d_1_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_56 = _T_6928 ? io_sc2mac_dat_mask_56 : in_rt_dat_mask_d_1_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_57 = _T_6928 ? io_sc2mac_dat_mask_57 : in_rt_dat_mask_d_1_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_58 = _T_6928 ? io_sc2mac_dat_mask_58 : in_rt_dat_mask_d_1_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_59 = _T_6928 ? io_sc2mac_dat_mask_59 : in_rt_dat_mask_d_1_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_60 = _T_6928 ? io_sc2mac_dat_mask_60 : in_rt_dat_mask_d_1_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_61 = _T_6928 ? io_sc2mac_dat_mask_61 : in_rt_dat_mask_d_1_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_62 = _T_6928 ? io_sc2mac_dat_mask_62 : in_rt_dat_mask_d_1_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_63 = _T_6928 ? io_sc2mac_dat_mask_63 : in_rt_dat_mask_d_1_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_64 = _T_6928 ? io_sc2mac_dat_mask_64 : in_rt_dat_mask_d_1_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_65 = _T_6928 ? io_sc2mac_dat_mask_65 : in_rt_dat_mask_d_1_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_66 = _T_6928 ? io_sc2mac_dat_mask_66 : in_rt_dat_mask_d_1_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_67 = _T_6928 ? io_sc2mac_dat_mask_67 : in_rt_dat_mask_d_1_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_68 = _T_6928 ? io_sc2mac_dat_mask_68 : in_rt_dat_mask_d_1_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_69 = _T_6928 ? io_sc2mac_dat_mask_69 : in_rt_dat_mask_d_1_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_70 = _T_6928 ? io_sc2mac_dat_mask_70 : in_rt_dat_mask_d_1_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_71 = _T_6928 ? io_sc2mac_dat_mask_71 : in_rt_dat_mask_d_1_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_72 = _T_6928 ? io_sc2mac_dat_mask_72 : in_rt_dat_mask_d_1_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_73 = _T_6928 ? io_sc2mac_dat_mask_73 : in_rt_dat_mask_d_1_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_74 = _T_6928 ? io_sc2mac_dat_mask_74 : in_rt_dat_mask_d_1_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_75 = _T_6928 ? io_sc2mac_dat_mask_75 : in_rt_dat_mask_d_1_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_76 = _T_6928 ? io_sc2mac_dat_mask_76 : in_rt_dat_mask_d_1_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_77 = _T_6928 ? io_sc2mac_dat_mask_77 : in_rt_dat_mask_d_1_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_78 = _T_6928 ? io_sc2mac_dat_mask_78 : in_rt_dat_mask_d_1_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_79 = _T_6928 ? io_sc2mac_dat_mask_79 : in_rt_dat_mask_d_1_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_80 = _T_6928 ? io_sc2mac_dat_mask_80 : in_rt_dat_mask_d_1_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_81 = _T_6928 ? io_sc2mac_dat_mask_81 : in_rt_dat_mask_d_1_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_82 = _T_6928 ? io_sc2mac_dat_mask_82 : in_rt_dat_mask_d_1_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_83 = _T_6928 ? io_sc2mac_dat_mask_83 : in_rt_dat_mask_d_1_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_84 = _T_6928 ? io_sc2mac_dat_mask_84 : in_rt_dat_mask_d_1_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_85 = _T_6928 ? io_sc2mac_dat_mask_85 : in_rt_dat_mask_d_1_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_86 = _T_6928 ? io_sc2mac_dat_mask_86 : in_rt_dat_mask_d_1_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_87 = _T_6928 ? io_sc2mac_dat_mask_87 : in_rt_dat_mask_d_1_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_88 = _T_6928 ? io_sc2mac_dat_mask_88 : in_rt_dat_mask_d_1_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_89 = _T_6928 ? io_sc2mac_dat_mask_89 : in_rt_dat_mask_d_1_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_90 = _T_6928 ? io_sc2mac_dat_mask_90 : in_rt_dat_mask_d_1_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_91 = _T_6928 ? io_sc2mac_dat_mask_91 : in_rt_dat_mask_d_1_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_92 = _T_6928 ? io_sc2mac_dat_mask_92 : in_rt_dat_mask_d_1_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_93 = _T_6928 ? io_sc2mac_dat_mask_93 : in_rt_dat_mask_d_1_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_94 = _T_6928 ? io_sc2mac_dat_mask_94 : in_rt_dat_mask_d_1_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_95 = _T_6928 ? io_sc2mac_dat_mask_95 : in_rt_dat_mask_d_1_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_96 = _T_6928 ? io_sc2mac_dat_mask_96 : in_rt_dat_mask_d_1_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_97 = _T_6928 ? io_sc2mac_dat_mask_97 : in_rt_dat_mask_d_1_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_98 = _T_6928 ? io_sc2mac_dat_mask_98 : in_rt_dat_mask_d_1_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_99 = _T_6928 ? io_sc2mac_dat_mask_99 : in_rt_dat_mask_d_1_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_100 = _T_6928 ? io_sc2mac_dat_mask_100 : in_rt_dat_mask_d_1_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_101 = _T_6928 ? io_sc2mac_dat_mask_101 : in_rt_dat_mask_d_1_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_102 = _T_6928 ? io_sc2mac_dat_mask_102 : in_rt_dat_mask_d_1_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_103 = _T_6928 ? io_sc2mac_dat_mask_103 : in_rt_dat_mask_d_1_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_104 = _T_6928 ? io_sc2mac_dat_mask_104 : in_rt_dat_mask_d_1_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_105 = _T_6928 ? io_sc2mac_dat_mask_105 : in_rt_dat_mask_d_1_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_106 = _T_6928 ? io_sc2mac_dat_mask_106 : in_rt_dat_mask_d_1_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_107 = _T_6928 ? io_sc2mac_dat_mask_107 : in_rt_dat_mask_d_1_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_108 = _T_6928 ? io_sc2mac_dat_mask_108 : in_rt_dat_mask_d_1_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_109 = _T_6928 ? io_sc2mac_dat_mask_109 : in_rt_dat_mask_d_1_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_110 = _T_6928 ? io_sc2mac_dat_mask_110 : in_rt_dat_mask_d_1_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_111 = _T_6928 ? io_sc2mac_dat_mask_111 : in_rt_dat_mask_d_1_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_112 = _T_6928 ? io_sc2mac_dat_mask_112 : in_rt_dat_mask_d_1_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_113 = _T_6928 ? io_sc2mac_dat_mask_113 : in_rt_dat_mask_d_1_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_114 = _T_6928 ? io_sc2mac_dat_mask_114 : in_rt_dat_mask_d_1_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_115 = _T_6928 ? io_sc2mac_dat_mask_115 : in_rt_dat_mask_d_1_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_116 = _T_6928 ? io_sc2mac_dat_mask_116 : in_rt_dat_mask_d_1_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_117 = _T_6928 ? io_sc2mac_dat_mask_117 : in_rt_dat_mask_d_1_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_118 = _T_6928 ? io_sc2mac_dat_mask_118 : in_rt_dat_mask_d_1_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_119 = _T_6928 ? io_sc2mac_dat_mask_119 : in_rt_dat_mask_d_1_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_120 = _T_6928 ? io_sc2mac_dat_mask_120 : in_rt_dat_mask_d_1_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_121 = _T_6928 ? io_sc2mac_dat_mask_121 : in_rt_dat_mask_d_1_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_122 = _T_6928 ? io_sc2mac_dat_mask_122 : in_rt_dat_mask_d_1_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_123 = _T_6928 ? io_sc2mac_dat_mask_123 : in_rt_dat_mask_d_1_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_124 = _T_6928 ? io_sc2mac_dat_mask_124 : in_rt_dat_mask_d_1_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_125 = _T_6928 ? io_sc2mac_dat_mask_125 : in_rt_dat_mask_d_1_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_126 = _T_6928 ? io_sc2mac_dat_mask_126 : in_rt_dat_mask_d_1_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_127 = _T_6928 ? io_sc2mac_dat_mask_127 : in_rt_dat_mask_d_1_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_128 = _T_6928 ? io_sc2mac_dat_pd : in_rt_dat_pd_d_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _T_6929 = io_sc2mac_wt_pvld | in_rt_wt_pvld_d_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:32]
  assign _GEN_129 = _T_6929 ? io_sc2mac_wt_mask_0 : in_rt_wt_mask_d_1_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_130 = _T_6929 ? io_sc2mac_wt_mask_1 : in_rt_wt_mask_d_1_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_131 = _T_6929 ? io_sc2mac_wt_mask_2 : in_rt_wt_mask_d_1_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_132 = _T_6929 ? io_sc2mac_wt_mask_3 : in_rt_wt_mask_d_1_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_133 = _T_6929 ? io_sc2mac_wt_mask_4 : in_rt_wt_mask_d_1_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_134 = _T_6929 ? io_sc2mac_wt_mask_5 : in_rt_wt_mask_d_1_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_135 = _T_6929 ? io_sc2mac_wt_mask_6 : in_rt_wt_mask_d_1_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_136 = _T_6929 ? io_sc2mac_wt_mask_7 : in_rt_wt_mask_d_1_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_137 = _T_6929 ? io_sc2mac_wt_mask_8 : in_rt_wt_mask_d_1_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_138 = _T_6929 ? io_sc2mac_wt_mask_9 : in_rt_wt_mask_d_1_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_139 = _T_6929 ? io_sc2mac_wt_mask_10 : in_rt_wt_mask_d_1_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_140 = _T_6929 ? io_sc2mac_wt_mask_11 : in_rt_wt_mask_d_1_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_141 = _T_6929 ? io_sc2mac_wt_mask_12 : in_rt_wt_mask_d_1_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_142 = _T_6929 ? io_sc2mac_wt_mask_13 : in_rt_wt_mask_d_1_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_143 = _T_6929 ? io_sc2mac_wt_mask_14 : in_rt_wt_mask_d_1_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_144 = _T_6929 ? io_sc2mac_wt_mask_15 : in_rt_wt_mask_d_1_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_145 = _T_6929 ? io_sc2mac_wt_mask_16 : in_rt_wt_mask_d_1_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_146 = _T_6929 ? io_sc2mac_wt_mask_17 : in_rt_wt_mask_d_1_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_147 = _T_6929 ? io_sc2mac_wt_mask_18 : in_rt_wt_mask_d_1_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_148 = _T_6929 ? io_sc2mac_wt_mask_19 : in_rt_wt_mask_d_1_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_149 = _T_6929 ? io_sc2mac_wt_mask_20 : in_rt_wt_mask_d_1_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_150 = _T_6929 ? io_sc2mac_wt_mask_21 : in_rt_wt_mask_d_1_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_151 = _T_6929 ? io_sc2mac_wt_mask_22 : in_rt_wt_mask_d_1_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_152 = _T_6929 ? io_sc2mac_wt_mask_23 : in_rt_wt_mask_d_1_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_153 = _T_6929 ? io_sc2mac_wt_mask_24 : in_rt_wt_mask_d_1_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_154 = _T_6929 ? io_sc2mac_wt_mask_25 : in_rt_wt_mask_d_1_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_155 = _T_6929 ? io_sc2mac_wt_mask_26 : in_rt_wt_mask_d_1_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_156 = _T_6929 ? io_sc2mac_wt_mask_27 : in_rt_wt_mask_d_1_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_157 = _T_6929 ? io_sc2mac_wt_mask_28 : in_rt_wt_mask_d_1_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_158 = _T_6929 ? io_sc2mac_wt_mask_29 : in_rt_wt_mask_d_1_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_159 = _T_6929 ? io_sc2mac_wt_mask_30 : in_rt_wt_mask_d_1_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_160 = _T_6929 ? io_sc2mac_wt_mask_31 : in_rt_wt_mask_d_1_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_161 = _T_6929 ? io_sc2mac_wt_mask_32 : in_rt_wt_mask_d_1_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_162 = _T_6929 ? io_sc2mac_wt_mask_33 : in_rt_wt_mask_d_1_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_163 = _T_6929 ? io_sc2mac_wt_mask_34 : in_rt_wt_mask_d_1_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_164 = _T_6929 ? io_sc2mac_wt_mask_35 : in_rt_wt_mask_d_1_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_165 = _T_6929 ? io_sc2mac_wt_mask_36 : in_rt_wt_mask_d_1_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_166 = _T_6929 ? io_sc2mac_wt_mask_37 : in_rt_wt_mask_d_1_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_167 = _T_6929 ? io_sc2mac_wt_mask_38 : in_rt_wt_mask_d_1_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_168 = _T_6929 ? io_sc2mac_wt_mask_39 : in_rt_wt_mask_d_1_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_169 = _T_6929 ? io_sc2mac_wt_mask_40 : in_rt_wt_mask_d_1_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_170 = _T_6929 ? io_sc2mac_wt_mask_41 : in_rt_wt_mask_d_1_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_171 = _T_6929 ? io_sc2mac_wt_mask_42 : in_rt_wt_mask_d_1_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_172 = _T_6929 ? io_sc2mac_wt_mask_43 : in_rt_wt_mask_d_1_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_173 = _T_6929 ? io_sc2mac_wt_mask_44 : in_rt_wt_mask_d_1_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_174 = _T_6929 ? io_sc2mac_wt_mask_45 : in_rt_wt_mask_d_1_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_175 = _T_6929 ? io_sc2mac_wt_mask_46 : in_rt_wt_mask_d_1_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_176 = _T_6929 ? io_sc2mac_wt_mask_47 : in_rt_wt_mask_d_1_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_177 = _T_6929 ? io_sc2mac_wt_mask_48 : in_rt_wt_mask_d_1_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_178 = _T_6929 ? io_sc2mac_wt_mask_49 : in_rt_wt_mask_d_1_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_179 = _T_6929 ? io_sc2mac_wt_mask_50 : in_rt_wt_mask_d_1_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_180 = _T_6929 ? io_sc2mac_wt_mask_51 : in_rt_wt_mask_d_1_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_181 = _T_6929 ? io_sc2mac_wt_mask_52 : in_rt_wt_mask_d_1_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_182 = _T_6929 ? io_sc2mac_wt_mask_53 : in_rt_wt_mask_d_1_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_183 = _T_6929 ? io_sc2mac_wt_mask_54 : in_rt_wt_mask_d_1_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_184 = _T_6929 ? io_sc2mac_wt_mask_55 : in_rt_wt_mask_d_1_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_185 = _T_6929 ? io_sc2mac_wt_mask_56 : in_rt_wt_mask_d_1_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_186 = _T_6929 ? io_sc2mac_wt_mask_57 : in_rt_wt_mask_d_1_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_187 = _T_6929 ? io_sc2mac_wt_mask_58 : in_rt_wt_mask_d_1_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_188 = _T_6929 ? io_sc2mac_wt_mask_59 : in_rt_wt_mask_d_1_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_189 = _T_6929 ? io_sc2mac_wt_mask_60 : in_rt_wt_mask_d_1_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_190 = _T_6929 ? io_sc2mac_wt_mask_61 : in_rt_wt_mask_d_1_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_191 = _T_6929 ? io_sc2mac_wt_mask_62 : in_rt_wt_mask_d_1_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_192 = _T_6929 ? io_sc2mac_wt_mask_63 : in_rt_wt_mask_d_1_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_193 = _T_6929 ? io_sc2mac_wt_mask_64 : in_rt_wt_mask_d_1_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_194 = _T_6929 ? io_sc2mac_wt_mask_65 : in_rt_wt_mask_d_1_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_195 = _T_6929 ? io_sc2mac_wt_mask_66 : in_rt_wt_mask_d_1_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_196 = _T_6929 ? io_sc2mac_wt_mask_67 : in_rt_wt_mask_d_1_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_197 = _T_6929 ? io_sc2mac_wt_mask_68 : in_rt_wt_mask_d_1_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_198 = _T_6929 ? io_sc2mac_wt_mask_69 : in_rt_wt_mask_d_1_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_199 = _T_6929 ? io_sc2mac_wt_mask_70 : in_rt_wt_mask_d_1_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_200 = _T_6929 ? io_sc2mac_wt_mask_71 : in_rt_wt_mask_d_1_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_201 = _T_6929 ? io_sc2mac_wt_mask_72 : in_rt_wt_mask_d_1_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_202 = _T_6929 ? io_sc2mac_wt_mask_73 : in_rt_wt_mask_d_1_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_203 = _T_6929 ? io_sc2mac_wt_mask_74 : in_rt_wt_mask_d_1_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_204 = _T_6929 ? io_sc2mac_wt_mask_75 : in_rt_wt_mask_d_1_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_205 = _T_6929 ? io_sc2mac_wt_mask_76 : in_rt_wt_mask_d_1_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_206 = _T_6929 ? io_sc2mac_wt_mask_77 : in_rt_wt_mask_d_1_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_207 = _T_6929 ? io_sc2mac_wt_mask_78 : in_rt_wt_mask_d_1_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_208 = _T_6929 ? io_sc2mac_wt_mask_79 : in_rt_wt_mask_d_1_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_209 = _T_6929 ? io_sc2mac_wt_mask_80 : in_rt_wt_mask_d_1_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_210 = _T_6929 ? io_sc2mac_wt_mask_81 : in_rt_wt_mask_d_1_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_211 = _T_6929 ? io_sc2mac_wt_mask_82 : in_rt_wt_mask_d_1_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_212 = _T_6929 ? io_sc2mac_wt_mask_83 : in_rt_wt_mask_d_1_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_213 = _T_6929 ? io_sc2mac_wt_mask_84 : in_rt_wt_mask_d_1_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_214 = _T_6929 ? io_sc2mac_wt_mask_85 : in_rt_wt_mask_d_1_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_215 = _T_6929 ? io_sc2mac_wt_mask_86 : in_rt_wt_mask_d_1_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_216 = _T_6929 ? io_sc2mac_wt_mask_87 : in_rt_wt_mask_d_1_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_217 = _T_6929 ? io_sc2mac_wt_mask_88 : in_rt_wt_mask_d_1_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_218 = _T_6929 ? io_sc2mac_wt_mask_89 : in_rt_wt_mask_d_1_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_219 = _T_6929 ? io_sc2mac_wt_mask_90 : in_rt_wt_mask_d_1_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_220 = _T_6929 ? io_sc2mac_wt_mask_91 : in_rt_wt_mask_d_1_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_221 = _T_6929 ? io_sc2mac_wt_mask_92 : in_rt_wt_mask_d_1_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_222 = _T_6929 ? io_sc2mac_wt_mask_93 : in_rt_wt_mask_d_1_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_223 = _T_6929 ? io_sc2mac_wt_mask_94 : in_rt_wt_mask_d_1_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_224 = _T_6929 ? io_sc2mac_wt_mask_95 : in_rt_wt_mask_d_1_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_225 = _T_6929 ? io_sc2mac_wt_mask_96 : in_rt_wt_mask_d_1_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_226 = _T_6929 ? io_sc2mac_wt_mask_97 : in_rt_wt_mask_d_1_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_227 = _T_6929 ? io_sc2mac_wt_mask_98 : in_rt_wt_mask_d_1_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_228 = _T_6929 ? io_sc2mac_wt_mask_99 : in_rt_wt_mask_d_1_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_229 = _T_6929 ? io_sc2mac_wt_mask_100 : in_rt_wt_mask_d_1_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_230 = _T_6929 ? io_sc2mac_wt_mask_101 : in_rt_wt_mask_d_1_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_231 = _T_6929 ? io_sc2mac_wt_mask_102 : in_rt_wt_mask_d_1_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_232 = _T_6929 ? io_sc2mac_wt_mask_103 : in_rt_wt_mask_d_1_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_233 = _T_6929 ? io_sc2mac_wt_mask_104 : in_rt_wt_mask_d_1_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_234 = _T_6929 ? io_sc2mac_wt_mask_105 : in_rt_wt_mask_d_1_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_235 = _T_6929 ? io_sc2mac_wt_mask_106 : in_rt_wt_mask_d_1_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_236 = _T_6929 ? io_sc2mac_wt_mask_107 : in_rt_wt_mask_d_1_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_237 = _T_6929 ? io_sc2mac_wt_mask_108 : in_rt_wt_mask_d_1_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_238 = _T_6929 ? io_sc2mac_wt_mask_109 : in_rt_wt_mask_d_1_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_239 = _T_6929 ? io_sc2mac_wt_mask_110 : in_rt_wt_mask_d_1_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_240 = _T_6929 ? io_sc2mac_wt_mask_111 : in_rt_wt_mask_d_1_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_241 = _T_6929 ? io_sc2mac_wt_mask_112 : in_rt_wt_mask_d_1_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_242 = _T_6929 ? io_sc2mac_wt_mask_113 : in_rt_wt_mask_d_1_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_243 = _T_6929 ? io_sc2mac_wt_mask_114 : in_rt_wt_mask_d_1_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_244 = _T_6929 ? io_sc2mac_wt_mask_115 : in_rt_wt_mask_d_1_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_245 = _T_6929 ? io_sc2mac_wt_mask_116 : in_rt_wt_mask_d_1_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_246 = _T_6929 ? io_sc2mac_wt_mask_117 : in_rt_wt_mask_d_1_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_247 = _T_6929 ? io_sc2mac_wt_mask_118 : in_rt_wt_mask_d_1_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_248 = _T_6929 ? io_sc2mac_wt_mask_119 : in_rt_wt_mask_d_1_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_249 = _T_6929 ? io_sc2mac_wt_mask_120 : in_rt_wt_mask_d_1_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_250 = _T_6929 ? io_sc2mac_wt_mask_121 : in_rt_wt_mask_d_1_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_251 = _T_6929 ? io_sc2mac_wt_mask_122 : in_rt_wt_mask_d_1_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_252 = _T_6929 ? io_sc2mac_wt_mask_123 : in_rt_wt_mask_d_1_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_253 = _T_6929 ? io_sc2mac_wt_mask_124 : in_rt_wt_mask_d_1_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_254 = _T_6929 ? io_sc2mac_wt_mask_125 : in_rt_wt_mask_d_1_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_255 = _T_6929 ? io_sc2mac_wt_mask_126 : in_rt_wt_mask_d_1_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_256 = _T_6929 ? io_sc2mac_wt_mask_127 : in_rt_wt_mask_d_1_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_257 = _T_6929 ? io_sc2mac_wt_sel_0 : in_rt_wt_sel_d_1_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _T_6930 = in_rt_dat_pvld_d_1 | in_rt_dat_pvld_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:33]
  assign _GEN_514 = _T_6930 ? in_rt_dat_mask_d_1_0 : in_rt_dat_mask_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_515 = _T_6930 ? in_rt_dat_mask_d_1_1 : in_rt_dat_mask_d_2_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_516 = _T_6930 ? in_rt_dat_mask_d_1_2 : in_rt_dat_mask_d_2_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_517 = _T_6930 ? in_rt_dat_mask_d_1_3 : in_rt_dat_mask_d_2_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_518 = _T_6930 ? in_rt_dat_mask_d_1_4 : in_rt_dat_mask_d_2_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_519 = _T_6930 ? in_rt_dat_mask_d_1_5 : in_rt_dat_mask_d_2_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_520 = _T_6930 ? in_rt_dat_mask_d_1_6 : in_rt_dat_mask_d_2_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_521 = _T_6930 ? in_rt_dat_mask_d_1_7 : in_rt_dat_mask_d_2_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_522 = _T_6930 ? in_rt_dat_mask_d_1_8 : in_rt_dat_mask_d_2_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_523 = _T_6930 ? in_rt_dat_mask_d_1_9 : in_rt_dat_mask_d_2_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_524 = _T_6930 ? in_rt_dat_mask_d_1_10 : in_rt_dat_mask_d_2_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_525 = _T_6930 ? in_rt_dat_mask_d_1_11 : in_rt_dat_mask_d_2_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_526 = _T_6930 ? in_rt_dat_mask_d_1_12 : in_rt_dat_mask_d_2_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_527 = _T_6930 ? in_rt_dat_mask_d_1_13 : in_rt_dat_mask_d_2_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_528 = _T_6930 ? in_rt_dat_mask_d_1_14 : in_rt_dat_mask_d_2_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_529 = _T_6930 ? in_rt_dat_mask_d_1_15 : in_rt_dat_mask_d_2_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_530 = _T_6930 ? in_rt_dat_mask_d_1_16 : in_rt_dat_mask_d_2_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_531 = _T_6930 ? in_rt_dat_mask_d_1_17 : in_rt_dat_mask_d_2_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_532 = _T_6930 ? in_rt_dat_mask_d_1_18 : in_rt_dat_mask_d_2_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_533 = _T_6930 ? in_rt_dat_mask_d_1_19 : in_rt_dat_mask_d_2_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_534 = _T_6930 ? in_rt_dat_mask_d_1_20 : in_rt_dat_mask_d_2_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_535 = _T_6930 ? in_rt_dat_mask_d_1_21 : in_rt_dat_mask_d_2_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_536 = _T_6930 ? in_rt_dat_mask_d_1_22 : in_rt_dat_mask_d_2_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_537 = _T_6930 ? in_rt_dat_mask_d_1_23 : in_rt_dat_mask_d_2_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_538 = _T_6930 ? in_rt_dat_mask_d_1_24 : in_rt_dat_mask_d_2_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_539 = _T_6930 ? in_rt_dat_mask_d_1_25 : in_rt_dat_mask_d_2_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_540 = _T_6930 ? in_rt_dat_mask_d_1_26 : in_rt_dat_mask_d_2_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_541 = _T_6930 ? in_rt_dat_mask_d_1_27 : in_rt_dat_mask_d_2_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_542 = _T_6930 ? in_rt_dat_mask_d_1_28 : in_rt_dat_mask_d_2_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_543 = _T_6930 ? in_rt_dat_mask_d_1_29 : in_rt_dat_mask_d_2_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_544 = _T_6930 ? in_rt_dat_mask_d_1_30 : in_rt_dat_mask_d_2_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_545 = _T_6930 ? in_rt_dat_mask_d_1_31 : in_rt_dat_mask_d_2_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_546 = _T_6930 ? in_rt_dat_mask_d_1_32 : in_rt_dat_mask_d_2_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_547 = _T_6930 ? in_rt_dat_mask_d_1_33 : in_rt_dat_mask_d_2_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_548 = _T_6930 ? in_rt_dat_mask_d_1_34 : in_rt_dat_mask_d_2_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_549 = _T_6930 ? in_rt_dat_mask_d_1_35 : in_rt_dat_mask_d_2_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_550 = _T_6930 ? in_rt_dat_mask_d_1_36 : in_rt_dat_mask_d_2_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_551 = _T_6930 ? in_rt_dat_mask_d_1_37 : in_rt_dat_mask_d_2_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_552 = _T_6930 ? in_rt_dat_mask_d_1_38 : in_rt_dat_mask_d_2_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_553 = _T_6930 ? in_rt_dat_mask_d_1_39 : in_rt_dat_mask_d_2_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_554 = _T_6930 ? in_rt_dat_mask_d_1_40 : in_rt_dat_mask_d_2_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_555 = _T_6930 ? in_rt_dat_mask_d_1_41 : in_rt_dat_mask_d_2_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_556 = _T_6930 ? in_rt_dat_mask_d_1_42 : in_rt_dat_mask_d_2_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_557 = _T_6930 ? in_rt_dat_mask_d_1_43 : in_rt_dat_mask_d_2_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_558 = _T_6930 ? in_rt_dat_mask_d_1_44 : in_rt_dat_mask_d_2_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_559 = _T_6930 ? in_rt_dat_mask_d_1_45 : in_rt_dat_mask_d_2_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_560 = _T_6930 ? in_rt_dat_mask_d_1_46 : in_rt_dat_mask_d_2_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_561 = _T_6930 ? in_rt_dat_mask_d_1_47 : in_rt_dat_mask_d_2_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_562 = _T_6930 ? in_rt_dat_mask_d_1_48 : in_rt_dat_mask_d_2_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_563 = _T_6930 ? in_rt_dat_mask_d_1_49 : in_rt_dat_mask_d_2_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_564 = _T_6930 ? in_rt_dat_mask_d_1_50 : in_rt_dat_mask_d_2_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_565 = _T_6930 ? in_rt_dat_mask_d_1_51 : in_rt_dat_mask_d_2_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_566 = _T_6930 ? in_rt_dat_mask_d_1_52 : in_rt_dat_mask_d_2_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_567 = _T_6930 ? in_rt_dat_mask_d_1_53 : in_rt_dat_mask_d_2_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_568 = _T_6930 ? in_rt_dat_mask_d_1_54 : in_rt_dat_mask_d_2_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_569 = _T_6930 ? in_rt_dat_mask_d_1_55 : in_rt_dat_mask_d_2_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_570 = _T_6930 ? in_rt_dat_mask_d_1_56 : in_rt_dat_mask_d_2_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_571 = _T_6930 ? in_rt_dat_mask_d_1_57 : in_rt_dat_mask_d_2_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_572 = _T_6930 ? in_rt_dat_mask_d_1_58 : in_rt_dat_mask_d_2_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_573 = _T_6930 ? in_rt_dat_mask_d_1_59 : in_rt_dat_mask_d_2_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_574 = _T_6930 ? in_rt_dat_mask_d_1_60 : in_rt_dat_mask_d_2_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_575 = _T_6930 ? in_rt_dat_mask_d_1_61 : in_rt_dat_mask_d_2_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_576 = _T_6930 ? in_rt_dat_mask_d_1_62 : in_rt_dat_mask_d_2_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_577 = _T_6930 ? in_rt_dat_mask_d_1_63 : in_rt_dat_mask_d_2_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_578 = _T_6930 ? in_rt_dat_mask_d_1_64 : in_rt_dat_mask_d_2_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_579 = _T_6930 ? in_rt_dat_mask_d_1_65 : in_rt_dat_mask_d_2_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_580 = _T_6930 ? in_rt_dat_mask_d_1_66 : in_rt_dat_mask_d_2_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_581 = _T_6930 ? in_rt_dat_mask_d_1_67 : in_rt_dat_mask_d_2_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_582 = _T_6930 ? in_rt_dat_mask_d_1_68 : in_rt_dat_mask_d_2_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_583 = _T_6930 ? in_rt_dat_mask_d_1_69 : in_rt_dat_mask_d_2_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_584 = _T_6930 ? in_rt_dat_mask_d_1_70 : in_rt_dat_mask_d_2_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_585 = _T_6930 ? in_rt_dat_mask_d_1_71 : in_rt_dat_mask_d_2_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_586 = _T_6930 ? in_rt_dat_mask_d_1_72 : in_rt_dat_mask_d_2_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_587 = _T_6930 ? in_rt_dat_mask_d_1_73 : in_rt_dat_mask_d_2_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_588 = _T_6930 ? in_rt_dat_mask_d_1_74 : in_rt_dat_mask_d_2_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_589 = _T_6930 ? in_rt_dat_mask_d_1_75 : in_rt_dat_mask_d_2_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_590 = _T_6930 ? in_rt_dat_mask_d_1_76 : in_rt_dat_mask_d_2_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_591 = _T_6930 ? in_rt_dat_mask_d_1_77 : in_rt_dat_mask_d_2_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_592 = _T_6930 ? in_rt_dat_mask_d_1_78 : in_rt_dat_mask_d_2_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_593 = _T_6930 ? in_rt_dat_mask_d_1_79 : in_rt_dat_mask_d_2_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_594 = _T_6930 ? in_rt_dat_mask_d_1_80 : in_rt_dat_mask_d_2_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_595 = _T_6930 ? in_rt_dat_mask_d_1_81 : in_rt_dat_mask_d_2_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_596 = _T_6930 ? in_rt_dat_mask_d_1_82 : in_rt_dat_mask_d_2_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_597 = _T_6930 ? in_rt_dat_mask_d_1_83 : in_rt_dat_mask_d_2_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_598 = _T_6930 ? in_rt_dat_mask_d_1_84 : in_rt_dat_mask_d_2_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_599 = _T_6930 ? in_rt_dat_mask_d_1_85 : in_rt_dat_mask_d_2_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_600 = _T_6930 ? in_rt_dat_mask_d_1_86 : in_rt_dat_mask_d_2_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_601 = _T_6930 ? in_rt_dat_mask_d_1_87 : in_rt_dat_mask_d_2_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_602 = _T_6930 ? in_rt_dat_mask_d_1_88 : in_rt_dat_mask_d_2_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_603 = _T_6930 ? in_rt_dat_mask_d_1_89 : in_rt_dat_mask_d_2_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_604 = _T_6930 ? in_rt_dat_mask_d_1_90 : in_rt_dat_mask_d_2_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_605 = _T_6930 ? in_rt_dat_mask_d_1_91 : in_rt_dat_mask_d_2_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_606 = _T_6930 ? in_rt_dat_mask_d_1_92 : in_rt_dat_mask_d_2_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_607 = _T_6930 ? in_rt_dat_mask_d_1_93 : in_rt_dat_mask_d_2_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_608 = _T_6930 ? in_rt_dat_mask_d_1_94 : in_rt_dat_mask_d_2_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_609 = _T_6930 ? in_rt_dat_mask_d_1_95 : in_rt_dat_mask_d_2_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_610 = _T_6930 ? in_rt_dat_mask_d_1_96 : in_rt_dat_mask_d_2_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_611 = _T_6930 ? in_rt_dat_mask_d_1_97 : in_rt_dat_mask_d_2_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_612 = _T_6930 ? in_rt_dat_mask_d_1_98 : in_rt_dat_mask_d_2_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_613 = _T_6930 ? in_rt_dat_mask_d_1_99 : in_rt_dat_mask_d_2_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_614 = _T_6930 ? in_rt_dat_mask_d_1_100 : in_rt_dat_mask_d_2_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_615 = _T_6930 ? in_rt_dat_mask_d_1_101 : in_rt_dat_mask_d_2_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_616 = _T_6930 ? in_rt_dat_mask_d_1_102 : in_rt_dat_mask_d_2_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_617 = _T_6930 ? in_rt_dat_mask_d_1_103 : in_rt_dat_mask_d_2_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_618 = _T_6930 ? in_rt_dat_mask_d_1_104 : in_rt_dat_mask_d_2_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_619 = _T_6930 ? in_rt_dat_mask_d_1_105 : in_rt_dat_mask_d_2_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_620 = _T_6930 ? in_rt_dat_mask_d_1_106 : in_rt_dat_mask_d_2_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_621 = _T_6930 ? in_rt_dat_mask_d_1_107 : in_rt_dat_mask_d_2_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_622 = _T_6930 ? in_rt_dat_mask_d_1_108 : in_rt_dat_mask_d_2_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_623 = _T_6930 ? in_rt_dat_mask_d_1_109 : in_rt_dat_mask_d_2_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_624 = _T_6930 ? in_rt_dat_mask_d_1_110 : in_rt_dat_mask_d_2_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_625 = _T_6930 ? in_rt_dat_mask_d_1_111 : in_rt_dat_mask_d_2_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_626 = _T_6930 ? in_rt_dat_mask_d_1_112 : in_rt_dat_mask_d_2_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_627 = _T_6930 ? in_rt_dat_mask_d_1_113 : in_rt_dat_mask_d_2_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_628 = _T_6930 ? in_rt_dat_mask_d_1_114 : in_rt_dat_mask_d_2_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_629 = _T_6930 ? in_rt_dat_mask_d_1_115 : in_rt_dat_mask_d_2_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_630 = _T_6930 ? in_rt_dat_mask_d_1_116 : in_rt_dat_mask_d_2_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_631 = _T_6930 ? in_rt_dat_mask_d_1_117 : in_rt_dat_mask_d_2_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_632 = _T_6930 ? in_rt_dat_mask_d_1_118 : in_rt_dat_mask_d_2_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_633 = _T_6930 ? in_rt_dat_mask_d_1_119 : in_rt_dat_mask_d_2_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_634 = _T_6930 ? in_rt_dat_mask_d_1_120 : in_rt_dat_mask_d_2_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_635 = _T_6930 ? in_rt_dat_mask_d_1_121 : in_rt_dat_mask_d_2_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_636 = _T_6930 ? in_rt_dat_mask_d_1_122 : in_rt_dat_mask_d_2_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_637 = _T_6930 ? in_rt_dat_mask_d_1_123 : in_rt_dat_mask_d_2_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_638 = _T_6930 ? in_rt_dat_mask_d_1_124 : in_rt_dat_mask_d_2_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_639 = _T_6930 ? in_rt_dat_mask_d_1_125 : in_rt_dat_mask_d_2_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_640 = _T_6930 ? in_rt_dat_mask_d_1_126 : in_rt_dat_mask_d_2_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_641 = _T_6930 ? in_rt_dat_mask_d_1_127 : in_rt_dat_mask_d_2_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _GEN_642 = _T_6930 ? in_rt_dat_pd_d_1 : in_rt_dat_pd_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 92:56]
  assign _T_6931 = in_rt_wt_pvld_d_1 | in_rt_wt_pvld_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:32]
  assign _GEN_643 = _T_6931 ? in_rt_wt_mask_d_1_0 : in_rt_wt_mask_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_644 = _T_6931 ? in_rt_wt_mask_d_1_1 : in_rt_wt_mask_d_2_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_645 = _T_6931 ? in_rt_wt_mask_d_1_2 : in_rt_wt_mask_d_2_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_646 = _T_6931 ? in_rt_wt_mask_d_1_3 : in_rt_wt_mask_d_2_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_647 = _T_6931 ? in_rt_wt_mask_d_1_4 : in_rt_wt_mask_d_2_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_648 = _T_6931 ? in_rt_wt_mask_d_1_5 : in_rt_wt_mask_d_2_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_649 = _T_6931 ? in_rt_wt_mask_d_1_6 : in_rt_wt_mask_d_2_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_650 = _T_6931 ? in_rt_wt_mask_d_1_7 : in_rt_wt_mask_d_2_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_651 = _T_6931 ? in_rt_wt_mask_d_1_8 : in_rt_wt_mask_d_2_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_652 = _T_6931 ? in_rt_wt_mask_d_1_9 : in_rt_wt_mask_d_2_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_653 = _T_6931 ? in_rt_wt_mask_d_1_10 : in_rt_wt_mask_d_2_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_654 = _T_6931 ? in_rt_wt_mask_d_1_11 : in_rt_wt_mask_d_2_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_655 = _T_6931 ? in_rt_wt_mask_d_1_12 : in_rt_wt_mask_d_2_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_656 = _T_6931 ? in_rt_wt_mask_d_1_13 : in_rt_wt_mask_d_2_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_657 = _T_6931 ? in_rt_wt_mask_d_1_14 : in_rt_wt_mask_d_2_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_658 = _T_6931 ? in_rt_wt_mask_d_1_15 : in_rt_wt_mask_d_2_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_659 = _T_6931 ? in_rt_wt_mask_d_1_16 : in_rt_wt_mask_d_2_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_660 = _T_6931 ? in_rt_wt_mask_d_1_17 : in_rt_wt_mask_d_2_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_661 = _T_6931 ? in_rt_wt_mask_d_1_18 : in_rt_wt_mask_d_2_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_662 = _T_6931 ? in_rt_wt_mask_d_1_19 : in_rt_wt_mask_d_2_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_663 = _T_6931 ? in_rt_wt_mask_d_1_20 : in_rt_wt_mask_d_2_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_664 = _T_6931 ? in_rt_wt_mask_d_1_21 : in_rt_wt_mask_d_2_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_665 = _T_6931 ? in_rt_wt_mask_d_1_22 : in_rt_wt_mask_d_2_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_666 = _T_6931 ? in_rt_wt_mask_d_1_23 : in_rt_wt_mask_d_2_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_667 = _T_6931 ? in_rt_wt_mask_d_1_24 : in_rt_wt_mask_d_2_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_668 = _T_6931 ? in_rt_wt_mask_d_1_25 : in_rt_wt_mask_d_2_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_669 = _T_6931 ? in_rt_wt_mask_d_1_26 : in_rt_wt_mask_d_2_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_670 = _T_6931 ? in_rt_wt_mask_d_1_27 : in_rt_wt_mask_d_2_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_671 = _T_6931 ? in_rt_wt_mask_d_1_28 : in_rt_wt_mask_d_2_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_672 = _T_6931 ? in_rt_wt_mask_d_1_29 : in_rt_wt_mask_d_2_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_673 = _T_6931 ? in_rt_wt_mask_d_1_30 : in_rt_wt_mask_d_2_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_674 = _T_6931 ? in_rt_wt_mask_d_1_31 : in_rt_wt_mask_d_2_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_675 = _T_6931 ? in_rt_wt_mask_d_1_32 : in_rt_wt_mask_d_2_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_676 = _T_6931 ? in_rt_wt_mask_d_1_33 : in_rt_wt_mask_d_2_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_677 = _T_6931 ? in_rt_wt_mask_d_1_34 : in_rt_wt_mask_d_2_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_678 = _T_6931 ? in_rt_wt_mask_d_1_35 : in_rt_wt_mask_d_2_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_679 = _T_6931 ? in_rt_wt_mask_d_1_36 : in_rt_wt_mask_d_2_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_680 = _T_6931 ? in_rt_wt_mask_d_1_37 : in_rt_wt_mask_d_2_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_681 = _T_6931 ? in_rt_wt_mask_d_1_38 : in_rt_wt_mask_d_2_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_682 = _T_6931 ? in_rt_wt_mask_d_1_39 : in_rt_wt_mask_d_2_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_683 = _T_6931 ? in_rt_wt_mask_d_1_40 : in_rt_wt_mask_d_2_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_684 = _T_6931 ? in_rt_wt_mask_d_1_41 : in_rt_wt_mask_d_2_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_685 = _T_6931 ? in_rt_wt_mask_d_1_42 : in_rt_wt_mask_d_2_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_686 = _T_6931 ? in_rt_wt_mask_d_1_43 : in_rt_wt_mask_d_2_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_687 = _T_6931 ? in_rt_wt_mask_d_1_44 : in_rt_wt_mask_d_2_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_688 = _T_6931 ? in_rt_wt_mask_d_1_45 : in_rt_wt_mask_d_2_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_689 = _T_6931 ? in_rt_wt_mask_d_1_46 : in_rt_wt_mask_d_2_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_690 = _T_6931 ? in_rt_wt_mask_d_1_47 : in_rt_wt_mask_d_2_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_691 = _T_6931 ? in_rt_wt_mask_d_1_48 : in_rt_wt_mask_d_2_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_692 = _T_6931 ? in_rt_wt_mask_d_1_49 : in_rt_wt_mask_d_2_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_693 = _T_6931 ? in_rt_wt_mask_d_1_50 : in_rt_wt_mask_d_2_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_694 = _T_6931 ? in_rt_wt_mask_d_1_51 : in_rt_wt_mask_d_2_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_695 = _T_6931 ? in_rt_wt_mask_d_1_52 : in_rt_wt_mask_d_2_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_696 = _T_6931 ? in_rt_wt_mask_d_1_53 : in_rt_wt_mask_d_2_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_697 = _T_6931 ? in_rt_wt_mask_d_1_54 : in_rt_wt_mask_d_2_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_698 = _T_6931 ? in_rt_wt_mask_d_1_55 : in_rt_wt_mask_d_2_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_699 = _T_6931 ? in_rt_wt_mask_d_1_56 : in_rt_wt_mask_d_2_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_700 = _T_6931 ? in_rt_wt_mask_d_1_57 : in_rt_wt_mask_d_2_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_701 = _T_6931 ? in_rt_wt_mask_d_1_58 : in_rt_wt_mask_d_2_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_702 = _T_6931 ? in_rt_wt_mask_d_1_59 : in_rt_wt_mask_d_2_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_703 = _T_6931 ? in_rt_wt_mask_d_1_60 : in_rt_wt_mask_d_2_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_704 = _T_6931 ? in_rt_wt_mask_d_1_61 : in_rt_wt_mask_d_2_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_705 = _T_6931 ? in_rt_wt_mask_d_1_62 : in_rt_wt_mask_d_2_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_706 = _T_6931 ? in_rt_wt_mask_d_1_63 : in_rt_wt_mask_d_2_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_707 = _T_6931 ? in_rt_wt_mask_d_1_64 : in_rt_wt_mask_d_2_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_708 = _T_6931 ? in_rt_wt_mask_d_1_65 : in_rt_wt_mask_d_2_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_709 = _T_6931 ? in_rt_wt_mask_d_1_66 : in_rt_wt_mask_d_2_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_710 = _T_6931 ? in_rt_wt_mask_d_1_67 : in_rt_wt_mask_d_2_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_711 = _T_6931 ? in_rt_wt_mask_d_1_68 : in_rt_wt_mask_d_2_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_712 = _T_6931 ? in_rt_wt_mask_d_1_69 : in_rt_wt_mask_d_2_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_713 = _T_6931 ? in_rt_wt_mask_d_1_70 : in_rt_wt_mask_d_2_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_714 = _T_6931 ? in_rt_wt_mask_d_1_71 : in_rt_wt_mask_d_2_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_715 = _T_6931 ? in_rt_wt_mask_d_1_72 : in_rt_wt_mask_d_2_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_716 = _T_6931 ? in_rt_wt_mask_d_1_73 : in_rt_wt_mask_d_2_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_717 = _T_6931 ? in_rt_wt_mask_d_1_74 : in_rt_wt_mask_d_2_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_718 = _T_6931 ? in_rt_wt_mask_d_1_75 : in_rt_wt_mask_d_2_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_719 = _T_6931 ? in_rt_wt_mask_d_1_76 : in_rt_wt_mask_d_2_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_720 = _T_6931 ? in_rt_wt_mask_d_1_77 : in_rt_wt_mask_d_2_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_721 = _T_6931 ? in_rt_wt_mask_d_1_78 : in_rt_wt_mask_d_2_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_722 = _T_6931 ? in_rt_wt_mask_d_1_79 : in_rt_wt_mask_d_2_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_723 = _T_6931 ? in_rt_wt_mask_d_1_80 : in_rt_wt_mask_d_2_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_724 = _T_6931 ? in_rt_wt_mask_d_1_81 : in_rt_wt_mask_d_2_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_725 = _T_6931 ? in_rt_wt_mask_d_1_82 : in_rt_wt_mask_d_2_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_726 = _T_6931 ? in_rt_wt_mask_d_1_83 : in_rt_wt_mask_d_2_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_727 = _T_6931 ? in_rt_wt_mask_d_1_84 : in_rt_wt_mask_d_2_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_728 = _T_6931 ? in_rt_wt_mask_d_1_85 : in_rt_wt_mask_d_2_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_729 = _T_6931 ? in_rt_wt_mask_d_1_86 : in_rt_wt_mask_d_2_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_730 = _T_6931 ? in_rt_wt_mask_d_1_87 : in_rt_wt_mask_d_2_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_731 = _T_6931 ? in_rt_wt_mask_d_1_88 : in_rt_wt_mask_d_2_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_732 = _T_6931 ? in_rt_wt_mask_d_1_89 : in_rt_wt_mask_d_2_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_733 = _T_6931 ? in_rt_wt_mask_d_1_90 : in_rt_wt_mask_d_2_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_734 = _T_6931 ? in_rt_wt_mask_d_1_91 : in_rt_wt_mask_d_2_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_735 = _T_6931 ? in_rt_wt_mask_d_1_92 : in_rt_wt_mask_d_2_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_736 = _T_6931 ? in_rt_wt_mask_d_1_93 : in_rt_wt_mask_d_2_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_737 = _T_6931 ? in_rt_wt_mask_d_1_94 : in_rt_wt_mask_d_2_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_738 = _T_6931 ? in_rt_wt_mask_d_1_95 : in_rt_wt_mask_d_2_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_739 = _T_6931 ? in_rt_wt_mask_d_1_96 : in_rt_wt_mask_d_2_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_740 = _T_6931 ? in_rt_wt_mask_d_1_97 : in_rt_wt_mask_d_2_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_741 = _T_6931 ? in_rt_wt_mask_d_1_98 : in_rt_wt_mask_d_2_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_742 = _T_6931 ? in_rt_wt_mask_d_1_99 : in_rt_wt_mask_d_2_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_743 = _T_6931 ? in_rt_wt_mask_d_1_100 : in_rt_wt_mask_d_2_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_744 = _T_6931 ? in_rt_wt_mask_d_1_101 : in_rt_wt_mask_d_2_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_745 = _T_6931 ? in_rt_wt_mask_d_1_102 : in_rt_wt_mask_d_2_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_746 = _T_6931 ? in_rt_wt_mask_d_1_103 : in_rt_wt_mask_d_2_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_747 = _T_6931 ? in_rt_wt_mask_d_1_104 : in_rt_wt_mask_d_2_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_748 = _T_6931 ? in_rt_wt_mask_d_1_105 : in_rt_wt_mask_d_2_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_749 = _T_6931 ? in_rt_wt_mask_d_1_106 : in_rt_wt_mask_d_2_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_750 = _T_6931 ? in_rt_wt_mask_d_1_107 : in_rt_wt_mask_d_2_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_751 = _T_6931 ? in_rt_wt_mask_d_1_108 : in_rt_wt_mask_d_2_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_752 = _T_6931 ? in_rt_wt_mask_d_1_109 : in_rt_wt_mask_d_2_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_753 = _T_6931 ? in_rt_wt_mask_d_1_110 : in_rt_wt_mask_d_2_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_754 = _T_6931 ? in_rt_wt_mask_d_1_111 : in_rt_wt_mask_d_2_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_755 = _T_6931 ? in_rt_wt_mask_d_1_112 : in_rt_wt_mask_d_2_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_756 = _T_6931 ? in_rt_wt_mask_d_1_113 : in_rt_wt_mask_d_2_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_757 = _T_6931 ? in_rt_wt_mask_d_1_114 : in_rt_wt_mask_d_2_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_758 = _T_6931 ? in_rt_wt_mask_d_1_115 : in_rt_wt_mask_d_2_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_759 = _T_6931 ? in_rt_wt_mask_d_1_116 : in_rt_wt_mask_d_2_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_760 = _T_6931 ? in_rt_wt_mask_d_1_117 : in_rt_wt_mask_d_2_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_761 = _T_6931 ? in_rt_wt_mask_d_1_118 : in_rt_wt_mask_d_2_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_762 = _T_6931 ? in_rt_wt_mask_d_1_119 : in_rt_wt_mask_d_2_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_763 = _T_6931 ? in_rt_wt_mask_d_1_120 : in_rt_wt_mask_d_2_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_764 = _T_6931 ? in_rt_wt_mask_d_1_121 : in_rt_wt_mask_d_2_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_765 = _T_6931 ? in_rt_wt_mask_d_1_122 : in_rt_wt_mask_d_2_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_766 = _T_6931 ? in_rt_wt_mask_d_1_123 : in_rt_wt_mask_d_2_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_767 = _T_6931 ? in_rt_wt_mask_d_1_124 : in_rt_wt_mask_d_2_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_768 = _T_6931 ? in_rt_wt_mask_d_1_125 : in_rt_wt_mask_d_2_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_769 = _T_6931 ? in_rt_wt_mask_d_1_126 : in_rt_wt_mask_d_2_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_770 = _T_6931 ? in_rt_wt_mask_d_1_127 : in_rt_wt_mask_d_2_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign _GEN_771 = _T_6931 ? in_rt_wt_sel_d_1_0 : in_rt_wt_sel_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 98:54]
  assign io_in_dat_data_0 = in_rt_dat_data_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_1 = in_rt_dat_data_d_2_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_2 = in_rt_dat_data_d_2_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_3 = in_rt_dat_data_d_2_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_4 = in_rt_dat_data_d_2_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_5 = in_rt_dat_data_d_2_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_6 = in_rt_dat_data_d_2_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_7 = in_rt_dat_data_d_2_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_8 = in_rt_dat_data_d_2_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_9 = in_rt_dat_data_d_2_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_10 = in_rt_dat_data_d_2_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_11 = in_rt_dat_data_d_2_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_12 = in_rt_dat_data_d_2_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_13 = in_rt_dat_data_d_2_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_14 = in_rt_dat_data_d_2_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_15 = in_rt_dat_data_d_2_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_16 = in_rt_dat_data_d_2_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_17 = in_rt_dat_data_d_2_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_18 = in_rt_dat_data_d_2_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_19 = in_rt_dat_data_d_2_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_20 = in_rt_dat_data_d_2_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_21 = in_rt_dat_data_d_2_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_22 = in_rt_dat_data_d_2_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_23 = in_rt_dat_data_d_2_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_24 = in_rt_dat_data_d_2_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_25 = in_rt_dat_data_d_2_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_26 = in_rt_dat_data_d_2_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_27 = in_rt_dat_data_d_2_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_28 = in_rt_dat_data_d_2_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_29 = in_rt_dat_data_d_2_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_30 = in_rt_dat_data_d_2_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_31 = in_rt_dat_data_d_2_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_32 = in_rt_dat_data_d_2_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_33 = in_rt_dat_data_d_2_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_34 = in_rt_dat_data_d_2_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_35 = in_rt_dat_data_d_2_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_36 = in_rt_dat_data_d_2_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_37 = in_rt_dat_data_d_2_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_38 = in_rt_dat_data_d_2_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_39 = in_rt_dat_data_d_2_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_40 = in_rt_dat_data_d_2_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_41 = in_rt_dat_data_d_2_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_42 = in_rt_dat_data_d_2_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_43 = in_rt_dat_data_d_2_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_44 = in_rt_dat_data_d_2_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_45 = in_rt_dat_data_d_2_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_46 = in_rt_dat_data_d_2_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_47 = in_rt_dat_data_d_2_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_48 = in_rt_dat_data_d_2_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_49 = in_rt_dat_data_d_2_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_50 = in_rt_dat_data_d_2_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_51 = in_rt_dat_data_d_2_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_52 = in_rt_dat_data_d_2_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_53 = in_rt_dat_data_d_2_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_54 = in_rt_dat_data_d_2_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_55 = in_rt_dat_data_d_2_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_56 = in_rt_dat_data_d_2_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_57 = in_rt_dat_data_d_2_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_58 = in_rt_dat_data_d_2_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_59 = in_rt_dat_data_d_2_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_60 = in_rt_dat_data_d_2_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_61 = in_rt_dat_data_d_2_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_62 = in_rt_dat_data_d_2_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_63 = in_rt_dat_data_d_2_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_64 = in_rt_dat_data_d_2_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_65 = in_rt_dat_data_d_2_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_66 = in_rt_dat_data_d_2_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_67 = in_rt_dat_data_d_2_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_68 = in_rt_dat_data_d_2_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_69 = in_rt_dat_data_d_2_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_70 = in_rt_dat_data_d_2_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_71 = in_rt_dat_data_d_2_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_72 = in_rt_dat_data_d_2_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_73 = in_rt_dat_data_d_2_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_74 = in_rt_dat_data_d_2_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_75 = in_rt_dat_data_d_2_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_76 = in_rt_dat_data_d_2_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_77 = in_rt_dat_data_d_2_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_78 = in_rt_dat_data_d_2_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_79 = in_rt_dat_data_d_2_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_80 = in_rt_dat_data_d_2_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_81 = in_rt_dat_data_d_2_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_82 = in_rt_dat_data_d_2_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_83 = in_rt_dat_data_d_2_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_84 = in_rt_dat_data_d_2_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_85 = in_rt_dat_data_d_2_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_86 = in_rt_dat_data_d_2_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_87 = in_rt_dat_data_d_2_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_88 = in_rt_dat_data_d_2_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_89 = in_rt_dat_data_d_2_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_90 = in_rt_dat_data_d_2_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_91 = in_rt_dat_data_d_2_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_92 = in_rt_dat_data_d_2_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_93 = in_rt_dat_data_d_2_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_94 = in_rt_dat_data_d_2_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_95 = in_rt_dat_data_d_2_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_96 = in_rt_dat_data_d_2_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_97 = in_rt_dat_data_d_2_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_98 = in_rt_dat_data_d_2_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_99 = in_rt_dat_data_d_2_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_100 = in_rt_dat_data_d_2_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_101 = in_rt_dat_data_d_2_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_102 = in_rt_dat_data_d_2_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_103 = in_rt_dat_data_d_2_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_104 = in_rt_dat_data_d_2_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_105 = in_rt_dat_data_d_2_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_106 = in_rt_dat_data_d_2_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_107 = in_rt_dat_data_d_2_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_108 = in_rt_dat_data_d_2_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_109 = in_rt_dat_data_d_2_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_110 = in_rt_dat_data_d_2_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_111 = in_rt_dat_data_d_2_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_112 = in_rt_dat_data_d_2_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_113 = in_rt_dat_data_d_2_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_114 = in_rt_dat_data_d_2_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_115 = in_rt_dat_data_d_2_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_116 = in_rt_dat_data_d_2_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_117 = in_rt_dat_data_d_2_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_118 = in_rt_dat_data_d_2_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_119 = in_rt_dat_data_d_2_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_120 = in_rt_dat_data_d_2_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_121 = in_rt_dat_data_d_2_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_122 = in_rt_dat_data_d_2_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_123 = in_rt_dat_data_d_2_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_124 = in_rt_dat_data_d_2_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_125 = in_rt_dat_data_d_2_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_126 = in_rt_dat_data_d_2_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_data_127 = in_rt_dat_data_d_2_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 120:20]
  assign io_in_dat_mask_0 = in_rt_dat_mask_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_1 = in_rt_dat_mask_d_2_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_2 = in_rt_dat_mask_d_2_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_3 = in_rt_dat_mask_d_2_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_4 = in_rt_dat_mask_d_2_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_5 = in_rt_dat_mask_d_2_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_6 = in_rt_dat_mask_d_2_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_7 = in_rt_dat_mask_d_2_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_8 = in_rt_dat_mask_d_2_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_9 = in_rt_dat_mask_d_2_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_10 = in_rt_dat_mask_d_2_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_11 = in_rt_dat_mask_d_2_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_12 = in_rt_dat_mask_d_2_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_13 = in_rt_dat_mask_d_2_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_14 = in_rt_dat_mask_d_2_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_15 = in_rt_dat_mask_d_2_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_16 = in_rt_dat_mask_d_2_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_17 = in_rt_dat_mask_d_2_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_18 = in_rt_dat_mask_d_2_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_19 = in_rt_dat_mask_d_2_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_20 = in_rt_dat_mask_d_2_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_21 = in_rt_dat_mask_d_2_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_22 = in_rt_dat_mask_d_2_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_23 = in_rt_dat_mask_d_2_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_24 = in_rt_dat_mask_d_2_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_25 = in_rt_dat_mask_d_2_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_26 = in_rt_dat_mask_d_2_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_27 = in_rt_dat_mask_d_2_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_28 = in_rt_dat_mask_d_2_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_29 = in_rt_dat_mask_d_2_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_30 = in_rt_dat_mask_d_2_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_31 = in_rt_dat_mask_d_2_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_32 = in_rt_dat_mask_d_2_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_33 = in_rt_dat_mask_d_2_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_34 = in_rt_dat_mask_d_2_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_35 = in_rt_dat_mask_d_2_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_36 = in_rt_dat_mask_d_2_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_37 = in_rt_dat_mask_d_2_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_38 = in_rt_dat_mask_d_2_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_39 = in_rt_dat_mask_d_2_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_40 = in_rt_dat_mask_d_2_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_41 = in_rt_dat_mask_d_2_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_42 = in_rt_dat_mask_d_2_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_43 = in_rt_dat_mask_d_2_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_44 = in_rt_dat_mask_d_2_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_45 = in_rt_dat_mask_d_2_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_46 = in_rt_dat_mask_d_2_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_47 = in_rt_dat_mask_d_2_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_48 = in_rt_dat_mask_d_2_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_49 = in_rt_dat_mask_d_2_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_50 = in_rt_dat_mask_d_2_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_51 = in_rt_dat_mask_d_2_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_52 = in_rt_dat_mask_d_2_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_53 = in_rt_dat_mask_d_2_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_54 = in_rt_dat_mask_d_2_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_55 = in_rt_dat_mask_d_2_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_56 = in_rt_dat_mask_d_2_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_57 = in_rt_dat_mask_d_2_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_58 = in_rt_dat_mask_d_2_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_59 = in_rt_dat_mask_d_2_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_60 = in_rt_dat_mask_d_2_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_61 = in_rt_dat_mask_d_2_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_62 = in_rt_dat_mask_d_2_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_63 = in_rt_dat_mask_d_2_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_64 = in_rt_dat_mask_d_2_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_65 = in_rt_dat_mask_d_2_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_66 = in_rt_dat_mask_d_2_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_67 = in_rt_dat_mask_d_2_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_68 = in_rt_dat_mask_d_2_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_69 = in_rt_dat_mask_d_2_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_70 = in_rt_dat_mask_d_2_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_71 = in_rt_dat_mask_d_2_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_72 = in_rt_dat_mask_d_2_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_73 = in_rt_dat_mask_d_2_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_74 = in_rt_dat_mask_d_2_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_75 = in_rt_dat_mask_d_2_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_76 = in_rt_dat_mask_d_2_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_77 = in_rt_dat_mask_d_2_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_78 = in_rt_dat_mask_d_2_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_79 = in_rt_dat_mask_d_2_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_80 = in_rt_dat_mask_d_2_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_81 = in_rt_dat_mask_d_2_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_82 = in_rt_dat_mask_d_2_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_83 = in_rt_dat_mask_d_2_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_84 = in_rt_dat_mask_d_2_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_85 = in_rt_dat_mask_d_2_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_86 = in_rt_dat_mask_d_2_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_87 = in_rt_dat_mask_d_2_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_88 = in_rt_dat_mask_d_2_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_89 = in_rt_dat_mask_d_2_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_90 = in_rt_dat_mask_d_2_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_91 = in_rt_dat_mask_d_2_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_92 = in_rt_dat_mask_d_2_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_93 = in_rt_dat_mask_d_2_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_94 = in_rt_dat_mask_d_2_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_95 = in_rt_dat_mask_d_2_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_96 = in_rt_dat_mask_d_2_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_97 = in_rt_dat_mask_d_2_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_98 = in_rt_dat_mask_d_2_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_99 = in_rt_dat_mask_d_2_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_100 = in_rt_dat_mask_d_2_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_101 = in_rt_dat_mask_d_2_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_102 = in_rt_dat_mask_d_2_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_103 = in_rt_dat_mask_d_2_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_104 = in_rt_dat_mask_d_2_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_105 = in_rt_dat_mask_d_2_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_106 = in_rt_dat_mask_d_2_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_107 = in_rt_dat_mask_d_2_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_108 = in_rt_dat_mask_d_2_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_109 = in_rt_dat_mask_d_2_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_110 = in_rt_dat_mask_d_2_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_111 = in_rt_dat_mask_d_2_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_112 = in_rt_dat_mask_d_2_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_113 = in_rt_dat_mask_d_2_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_114 = in_rt_dat_mask_d_2_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_115 = in_rt_dat_mask_d_2_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_116 = in_rt_dat_mask_d_2_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_117 = in_rt_dat_mask_d_2_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_118 = in_rt_dat_mask_d_2_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_119 = in_rt_dat_mask_d_2_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_120 = in_rt_dat_mask_d_2_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_121 = in_rt_dat_mask_d_2_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_122 = in_rt_dat_mask_d_2_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_123 = in_rt_dat_mask_d_2_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_124 = in_rt_dat_mask_d_2_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_125 = in_rt_dat_mask_d_2_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_126 = in_rt_dat_mask_d_2_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_mask_127 = in_rt_dat_mask_d_2_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 115:20]
  assign io_in_dat_pd = in_rt_dat_pd_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 116:18]
  assign io_in_dat_pvld = in_rt_dat_pvld_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 114:20]
  assign io_in_dat_stripe_st = io_in_dat_pd[5]; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 123:25]
  assign io_in_dat_stripe_end = io_in_dat_pd[6]; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 124:26]
  assign io_in_wt_data_0 = in_rt_wt_data_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_1 = in_rt_wt_data_d_2_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_2 = in_rt_wt_data_d_2_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_3 = in_rt_wt_data_d_2_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_4 = in_rt_wt_data_d_2_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_5 = in_rt_wt_data_d_2_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_6 = in_rt_wt_data_d_2_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_7 = in_rt_wt_data_d_2_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_8 = in_rt_wt_data_d_2_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_9 = in_rt_wt_data_d_2_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_10 = in_rt_wt_data_d_2_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_11 = in_rt_wt_data_d_2_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_12 = in_rt_wt_data_d_2_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_13 = in_rt_wt_data_d_2_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_14 = in_rt_wt_data_d_2_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_15 = in_rt_wt_data_d_2_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_16 = in_rt_wt_data_d_2_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_17 = in_rt_wt_data_d_2_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_18 = in_rt_wt_data_d_2_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_19 = in_rt_wt_data_d_2_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_20 = in_rt_wt_data_d_2_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_21 = in_rt_wt_data_d_2_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_22 = in_rt_wt_data_d_2_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_23 = in_rt_wt_data_d_2_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_24 = in_rt_wt_data_d_2_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_25 = in_rt_wt_data_d_2_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_26 = in_rt_wt_data_d_2_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_27 = in_rt_wt_data_d_2_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_28 = in_rt_wt_data_d_2_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_29 = in_rt_wt_data_d_2_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_30 = in_rt_wt_data_d_2_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_31 = in_rt_wt_data_d_2_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_32 = in_rt_wt_data_d_2_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_33 = in_rt_wt_data_d_2_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_34 = in_rt_wt_data_d_2_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_35 = in_rt_wt_data_d_2_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_36 = in_rt_wt_data_d_2_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_37 = in_rt_wt_data_d_2_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_38 = in_rt_wt_data_d_2_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_39 = in_rt_wt_data_d_2_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_40 = in_rt_wt_data_d_2_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_41 = in_rt_wt_data_d_2_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_42 = in_rt_wt_data_d_2_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_43 = in_rt_wt_data_d_2_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_44 = in_rt_wt_data_d_2_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_45 = in_rt_wt_data_d_2_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_46 = in_rt_wt_data_d_2_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_47 = in_rt_wt_data_d_2_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_48 = in_rt_wt_data_d_2_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_49 = in_rt_wt_data_d_2_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_50 = in_rt_wt_data_d_2_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_51 = in_rt_wt_data_d_2_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_52 = in_rt_wt_data_d_2_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_53 = in_rt_wt_data_d_2_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_54 = in_rt_wt_data_d_2_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_55 = in_rt_wt_data_d_2_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_56 = in_rt_wt_data_d_2_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_57 = in_rt_wt_data_d_2_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_58 = in_rt_wt_data_d_2_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_59 = in_rt_wt_data_d_2_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_60 = in_rt_wt_data_d_2_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_61 = in_rt_wt_data_d_2_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_62 = in_rt_wt_data_d_2_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_63 = in_rt_wt_data_d_2_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_64 = in_rt_wt_data_d_2_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_65 = in_rt_wt_data_d_2_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_66 = in_rt_wt_data_d_2_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_67 = in_rt_wt_data_d_2_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_68 = in_rt_wt_data_d_2_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_69 = in_rt_wt_data_d_2_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_70 = in_rt_wt_data_d_2_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_71 = in_rt_wt_data_d_2_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_72 = in_rt_wt_data_d_2_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_73 = in_rt_wt_data_d_2_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_74 = in_rt_wt_data_d_2_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_75 = in_rt_wt_data_d_2_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_76 = in_rt_wt_data_d_2_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_77 = in_rt_wt_data_d_2_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_78 = in_rt_wt_data_d_2_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_79 = in_rt_wt_data_d_2_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_80 = in_rt_wt_data_d_2_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_81 = in_rt_wt_data_d_2_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_82 = in_rt_wt_data_d_2_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_83 = in_rt_wt_data_d_2_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_84 = in_rt_wt_data_d_2_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_85 = in_rt_wt_data_d_2_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_86 = in_rt_wt_data_d_2_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_87 = in_rt_wt_data_d_2_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_88 = in_rt_wt_data_d_2_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_89 = in_rt_wt_data_d_2_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_90 = in_rt_wt_data_d_2_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_91 = in_rt_wt_data_d_2_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_92 = in_rt_wt_data_d_2_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_93 = in_rt_wt_data_d_2_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_94 = in_rt_wt_data_d_2_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_95 = in_rt_wt_data_d_2_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_96 = in_rt_wt_data_d_2_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_97 = in_rt_wt_data_d_2_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_98 = in_rt_wt_data_d_2_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_99 = in_rt_wt_data_d_2_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_100 = in_rt_wt_data_d_2_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_101 = in_rt_wt_data_d_2_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_102 = in_rt_wt_data_d_2_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_103 = in_rt_wt_data_d_2_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_104 = in_rt_wt_data_d_2_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_105 = in_rt_wt_data_d_2_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_106 = in_rt_wt_data_d_2_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_107 = in_rt_wt_data_d_2_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_108 = in_rt_wt_data_d_2_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_109 = in_rt_wt_data_d_2_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_110 = in_rt_wt_data_d_2_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_111 = in_rt_wt_data_d_2_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_112 = in_rt_wt_data_d_2_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_113 = in_rt_wt_data_d_2_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_114 = in_rt_wt_data_d_2_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_115 = in_rt_wt_data_d_2_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_116 = in_rt_wt_data_d_2_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_117 = in_rt_wt_data_d_2_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_118 = in_rt_wt_data_d_2_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_119 = in_rt_wt_data_d_2_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_120 = in_rt_wt_data_d_2_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_121 = in_rt_wt_data_d_2_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_122 = in_rt_wt_data_d_2_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_123 = in_rt_wt_data_d_2_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_124 = in_rt_wt_data_d_2_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_125 = in_rt_wt_data_d_2_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_126 = in_rt_wt_data_d_2_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_data_127 = in_rt_wt_data_d_2_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 121:19]
  assign io_in_wt_mask_0 = in_rt_wt_mask_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_1 = in_rt_wt_mask_d_2_1; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_2 = in_rt_wt_mask_d_2_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_3 = in_rt_wt_mask_d_2_3; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_4 = in_rt_wt_mask_d_2_4; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_5 = in_rt_wt_mask_d_2_5; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_6 = in_rt_wt_mask_d_2_6; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_7 = in_rt_wt_mask_d_2_7; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_8 = in_rt_wt_mask_d_2_8; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_9 = in_rt_wt_mask_d_2_9; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_10 = in_rt_wt_mask_d_2_10; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_11 = in_rt_wt_mask_d_2_11; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_12 = in_rt_wt_mask_d_2_12; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_13 = in_rt_wt_mask_d_2_13; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_14 = in_rt_wt_mask_d_2_14; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_15 = in_rt_wt_mask_d_2_15; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_16 = in_rt_wt_mask_d_2_16; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_17 = in_rt_wt_mask_d_2_17; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_18 = in_rt_wt_mask_d_2_18; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_19 = in_rt_wt_mask_d_2_19; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_20 = in_rt_wt_mask_d_2_20; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_21 = in_rt_wt_mask_d_2_21; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_22 = in_rt_wt_mask_d_2_22; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_23 = in_rt_wt_mask_d_2_23; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_24 = in_rt_wt_mask_d_2_24; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_25 = in_rt_wt_mask_d_2_25; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_26 = in_rt_wt_mask_d_2_26; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_27 = in_rt_wt_mask_d_2_27; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_28 = in_rt_wt_mask_d_2_28; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_29 = in_rt_wt_mask_d_2_29; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_30 = in_rt_wt_mask_d_2_30; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_31 = in_rt_wt_mask_d_2_31; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_32 = in_rt_wt_mask_d_2_32; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_33 = in_rt_wt_mask_d_2_33; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_34 = in_rt_wt_mask_d_2_34; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_35 = in_rt_wt_mask_d_2_35; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_36 = in_rt_wt_mask_d_2_36; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_37 = in_rt_wt_mask_d_2_37; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_38 = in_rt_wt_mask_d_2_38; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_39 = in_rt_wt_mask_d_2_39; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_40 = in_rt_wt_mask_d_2_40; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_41 = in_rt_wt_mask_d_2_41; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_42 = in_rt_wt_mask_d_2_42; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_43 = in_rt_wt_mask_d_2_43; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_44 = in_rt_wt_mask_d_2_44; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_45 = in_rt_wt_mask_d_2_45; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_46 = in_rt_wt_mask_d_2_46; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_47 = in_rt_wt_mask_d_2_47; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_48 = in_rt_wt_mask_d_2_48; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_49 = in_rt_wt_mask_d_2_49; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_50 = in_rt_wt_mask_d_2_50; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_51 = in_rt_wt_mask_d_2_51; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_52 = in_rt_wt_mask_d_2_52; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_53 = in_rt_wt_mask_d_2_53; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_54 = in_rt_wt_mask_d_2_54; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_55 = in_rt_wt_mask_d_2_55; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_56 = in_rt_wt_mask_d_2_56; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_57 = in_rt_wt_mask_d_2_57; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_58 = in_rt_wt_mask_d_2_58; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_59 = in_rt_wt_mask_d_2_59; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_60 = in_rt_wt_mask_d_2_60; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_61 = in_rt_wt_mask_d_2_61; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_62 = in_rt_wt_mask_d_2_62; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_63 = in_rt_wt_mask_d_2_63; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_64 = in_rt_wt_mask_d_2_64; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_65 = in_rt_wt_mask_d_2_65; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_66 = in_rt_wt_mask_d_2_66; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_67 = in_rt_wt_mask_d_2_67; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_68 = in_rt_wt_mask_d_2_68; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_69 = in_rt_wt_mask_d_2_69; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_70 = in_rt_wt_mask_d_2_70; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_71 = in_rt_wt_mask_d_2_71; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_72 = in_rt_wt_mask_d_2_72; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_73 = in_rt_wt_mask_d_2_73; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_74 = in_rt_wt_mask_d_2_74; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_75 = in_rt_wt_mask_d_2_75; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_76 = in_rt_wt_mask_d_2_76; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_77 = in_rt_wt_mask_d_2_77; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_78 = in_rt_wt_mask_d_2_78; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_79 = in_rt_wt_mask_d_2_79; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_80 = in_rt_wt_mask_d_2_80; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_81 = in_rt_wt_mask_d_2_81; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_82 = in_rt_wt_mask_d_2_82; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_83 = in_rt_wt_mask_d_2_83; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_84 = in_rt_wt_mask_d_2_84; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_85 = in_rt_wt_mask_d_2_85; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_86 = in_rt_wt_mask_d_2_86; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_87 = in_rt_wt_mask_d_2_87; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_88 = in_rt_wt_mask_d_2_88; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_89 = in_rt_wt_mask_d_2_89; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_90 = in_rt_wt_mask_d_2_90; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_91 = in_rt_wt_mask_d_2_91; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_92 = in_rt_wt_mask_d_2_92; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_93 = in_rt_wt_mask_d_2_93; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_94 = in_rt_wt_mask_d_2_94; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_95 = in_rt_wt_mask_d_2_95; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_96 = in_rt_wt_mask_d_2_96; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_97 = in_rt_wt_mask_d_2_97; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_98 = in_rt_wt_mask_d_2_98; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_99 = in_rt_wt_mask_d_2_99; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_100 = in_rt_wt_mask_d_2_100; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_101 = in_rt_wt_mask_d_2_101; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_102 = in_rt_wt_mask_d_2_102; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_103 = in_rt_wt_mask_d_2_103; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_104 = in_rt_wt_mask_d_2_104; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_105 = in_rt_wt_mask_d_2_105; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_106 = in_rt_wt_mask_d_2_106; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_107 = in_rt_wt_mask_d_2_107; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_108 = in_rt_wt_mask_d_2_108; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_109 = in_rt_wt_mask_d_2_109; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_110 = in_rt_wt_mask_d_2_110; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_111 = in_rt_wt_mask_d_2_111; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_112 = in_rt_wt_mask_d_2_112; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_113 = in_rt_wt_mask_d_2_113; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_114 = in_rt_wt_mask_d_2_114; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_115 = in_rt_wt_mask_d_2_115; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_116 = in_rt_wt_mask_d_2_116; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_117 = in_rt_wt_mask_d_2_117; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_118 = in_rt_wt_mask_d_2_118; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_119 = in_rt_wt_mask_d_2_119; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_120 = in_rt_wt_mask_d_2_120; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_121 = in_rt_wt_mask_d_2_121; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_122 = in_rt_wt_mask_d_2_122; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_123 = in_rt_wt_mask_d_2_123; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_124 = in_rt_wt_mask_d_2_124; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_125 = in_rt_wt_mask_d_2_125; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_126 = in_rt_wt_mask_d_2_126; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_mask_127 = in_rt_wt_mask_d_2_127; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 118:19]
  assign io_in_wt_sel_0 = in_rt_wt_sel_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 119:18]
  assign io_in_wt_pvld = in_rt_wt_pvld_d_2; // @[NV_NVDLA_CMAC_CORE_rt_in.scala 117:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_rt_dat_data_d_1_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_rt_dat_data_d_1_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_rt_dat_data_d_1_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_rt_dat_data_d_1_3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_rt_dat_data_d_1_4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_rt_dat_data_d_1_5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  in_rt_dat_data_d_1_6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  in_rt_dat_data_d_1_7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  in_rt_dat_data_d_1_8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_rt_dat_data_d_1_9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_rt_dat_data_d_1_10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_rt_dat_data_d_1_11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_rt_dat_data_d_1_12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_rt_dat_data_d_1_13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_rt_dat_data_d_1_14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_rt_dat_data_d_1_15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_rt_dat_data_d_1_16 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_rt_dat_data_d_1_17 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_rt_dat_data_d_1_18 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_rt_dat_data_d_1_19 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_rt_dat_data_d_1_20 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_rt_dat_data_d_1_21 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_rt_dat_data_d_1_22 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_rt_dat_data_d_1_23 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_rt_dat_data_d_1_24 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_rt_dat_data_d_1_25 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  in_rt_dat_data_d_1_26 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  in_rt_dat_data_d_1_27 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  in_rt_dat_data_d_1_28 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  in_rt_dat_data_d_1_29 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  in_rt_dat_data_d_1_30 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  in_rt_dat_data_d_1_31 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  in_rt_dat_data_d_1_32 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  in_rt_dat_data_d_1_33 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  in_rt_dat_data_d_1_34 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  in_rt_dat_data_d_1_35 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  in_rt_dat_data_d_1_36 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  in_rt_dat_data_d_1_37 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  in_rt_dat_data_d_1_38 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  in_rt_dat_data_d_1_39 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  in_rt_dat_data_d_1_40 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  in_rt_dat_data_d_1_41 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  in_rt_dat_data_d_1_42 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  in_rt_dat_data_d_1_43 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  in_rt_dat_data_d_1_44 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  in_rt_dat_data_d_1_45 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  in_rt_dat_data_d_1_46 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  in_rt_dat_data_d_1_47 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  in_rt_dat_data_d_1_48 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  in_rt_dat_data_d_1_49 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  in_rt_dat_data_d_1_50 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  in_rt_dat_data_d_1_51 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  in_rt_dat_data_d_1_52 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  in_rt_dat_data_d_1_53 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  in_rt_dat_data_d_1_54 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  in_rt_dat_data_d_1_55 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  in_rt_dat_data_d_1_56 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  in_rt_dat_data_d_1_57 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  in_rt_dat_data_d_1_58 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  in_rt_dat_data_d_1_59 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  in_rt_dat_data_d_1_60 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  in_rt_dat_data_d_1_61 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  in_rt_dat_data_d_1_62 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  in_rt_dat_data_d_1_63 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  in_rt_dat_data_d_1_64 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  in_rt_dat_data_d_1_65 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  in_rt_dat_data_d_1_66 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  in_rt_dat_data_d_1_67 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  in_rt_dat_data_d_1_68 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  in_rt_dat_data_d_1_69 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  in_rt_dat_data_d_1_70 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  in_rt_dat_data_d_1_71 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  in_rt_dat_data_d_1_72 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  in_rt_dat_data_d_1_73 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  in_rt_dat_data_d_1_74 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  in_rt_dat_data_d_1_75 = _RAND_75[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  in_rt_dat_data_d_1_76 = _RAND_76[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  in_rt_dat_data_d_1_77 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  in_rt_dat_data_d_1_78 = _RAND_78[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  in_rt_dat_data_d_1_79 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  in_rt_dat_data_d_1_80 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  in_rt_dat_data_d_1_81 = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  in_rt_dat_data_d_1_82 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  in_rt_dat_data_d_1_83 = _RAND_83[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  in_rt_dat_data_d_1_84 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  in_rt_dat_data_d_1_85 = _RAND_85[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  in_rt_dat_data_d_1_86 = _RAND_86[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  in_rt_dat_data_d_1_87 = _RAND_87[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  in_rt_dat_data_d_1_88 = _RAND_88[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  in_rt_dat_data_d_1_89 = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  in_rt_dat_data_d_1_90 = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  in_rt_dat_data_d_1_91 = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  in_rt_dat_data_d_1_92 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  in_rt_dat_data_d_1_93 = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  in_rt_dat_data_d_1_94 = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  in_rt_dat_data_d_1_95 = _RAND_95[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  in_rt_dat_data_d_1_96 = _RAND_96[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  in_rt_dat_data_d_1_97 = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  in_rt_dat_data_d_1_98 = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  in_rt_dat_data_d_1_99 = _RAND_99[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  in_rt_dat_data_d_1_100 = _RAND_100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  in_rt_dat_data_d_1_101 = _RAND_101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  in_rt_dat_data_d_1_102 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  in_rt_dat_data_d_1_103 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  in_rt_dat_data_d_1_104 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  in_rt_dat_data_d_1_105 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  in_rt_dat_data_d_1_106 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  in_rt_dat_data_d_1_107 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  in_rt_dat_data_d_1_108 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  in_rt_dat_data_d_1_109 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  in_rt_dat_data_d_1_110 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  in_rt_dat_data_d_1_111 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  in_rt_dat_data_d_1_112 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  in_rt_dat_data_d_1_113 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  in_rt_dat_data_d_1_114 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  in_rt_dat_data_d_1_115 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  in_rt_dat_data_d_1_116 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  in_rt_dat_data_d_1_117 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  in_rt_dat_data_d_1_118 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  in_rt_dat_data_d_1_119 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  in_rt_dat_data_d_1_120 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  in_rt_dat_data_d_1_121 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  in_rt_dat_data_d_1_122 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  in_rt_dat_data_d_1_123 = _RAND_123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  in_rt_dat_data_d_1_124 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  in_rt_dat_data_d_1_125 = _RAND_125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  in_rt_dat_data_d_1_126 = _RAND_126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  in_rt_dat_data_d_1_127 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  in_rt_dat_data_d_2_0 = _RAND_128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  in_rt_dat_data_d_2_1 = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  in_rt_dat_data_d_2_2 = _RAND_130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  in_rt_dat_data_d_2_3 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  in_rt_dat_data_d_2_4 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  in_rt_dat_data_d_2_5 = _RAND_133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  in_rt_dat_data_d_2_6 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  in_rt_dat_data_d_2_7 = _RAND_135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  in_rt_dat_data_d_2_8 = _RAND_136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  in_rt_dat_data_d_2_9 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  in_rt_dat_data_d_2_10 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  in_rt_dat_data_d_2_11 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  in_rt_dat_data_d_2_12 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  in_rt_dat_data_d_2_13 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  in_rt_dat_data_d_2_14 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  in_rt_dat_data_d_2_15 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  in_rt_dat_data_d_2_16 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  in_rt_dat_data_d_2_17 = _RAND_145[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  in_rt_dat_data_d_2_18 = _RAND_146[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  in_rt_dat_data_d_2_19 = _RAND_147[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  in_rt_dat_data_d_2_20 = _RAND_148[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  in_rt_dat_data_d_2_21 = _RAND_149[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  in_rt_dat_data_d_2_22 = _RAND_150[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  in_rt_dat_data_d_2_23 = _RAND_151[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  in_rt_dat_data_d_2_24 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  in_rt_dat_data_d_2_25 = _RAND_153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  in_rt_dat_data_d_2_26 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  in_rt_dat_data_d_2_27 = _RAND_155[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  in_rt_dat_data_d_2_28 = _RAND_156[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  in_rt_dat_data_d_2_29 = _RAND_157[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  in_rt_dat_data_d_2_30 = _RAND_158[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  in_rt_dat_data_d_2_31 = _RAND_159[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  in_rt_dat_data_d_2_32 = _RAND_160[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  in_rt_dat_data_d_2_33 = _RAND_161[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  in_rt_dat_data_d_2_34 = _RAND_162[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  in_rt_dat_data_d_2_35 = _RAND_163[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  in_rt_dat_data_d_2_36 = _RAND_164[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  in_rt_dat_data_d_2_37 = _RAND_165[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  in_rt_dat_data_d_2_38 = _RAND_166[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  in_rt_dat_data_d_2_39 = _RAND_167[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  in_rt_dat_data_d_2_40 = _RAND_168[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  in_rt_dat_data_d_2_41 = _RAND_169[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  in_rt_dat_data_d_2_42 = _RAND_170[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  in_rt_dat_data_d_2_43 = _RAND_171[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  in_rt_dat_data_d_2_44 = _RAND_172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  in_rt_dat_data_d_2_45 = _RAND_173[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  in_rt_dat_data_d_2_46 = _RAND_174[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  in_rt_dat_data_d_2_47 = _RAND_175[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  in_rt_dat_data_d_2_48 = _RAND_176[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  in_rt_dat_data_d_2_49 = _RAND_177[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  in_rt_dat_data_d_2_50 = _RAND_178[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  in_rt_dat_data_d_2_51 = _RAND_179[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  in_rt_dat_data_d_2_52 = _RAND_180[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  in_rt_dat_data_d_2_53 = _RAND_181[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  in_rt_dat_data_d_2_54 = _RAND_182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  in_rt_dat_data_d_2_55 = _RAND_183[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  in_rt_dat_data_d_2_56 = _RAND_184[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  in_rt_dat_data_d_2_57 = _RAND_185[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  in_rt_dat_data_d_2_58 = _RAND_186[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  in_rt_dat_data_d_2_59 = _RAND_187[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  in_rt_dat_data_d_2_60 = _RAND_188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  in_rt_dat_data_d_2_61 = _RAND_189[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  in_rt_dat_data_d_2_62 = _RAND_190[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  in_rt_dat_data_d_2_63 = _RAND_191[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  in_rt_dat_data_d_2_64 = _RAND_192[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  in_rt_dat_data_d_2_65 = _RAND_193[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  in_rt_dat_data_d_2_66 = _RAND_194[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  in_rt_dat_data_d_2_67 = _RAND_195[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  in_rt_dat_data_d_2_68 = _RAND_196[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  in_rt_dat_data_d_2_69 = _RAND_197[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  in_rt_dat_data_d_2_70 = _RAND_198[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  in_rt_dat_data_d_2_71 = _RAND_199[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  in_rt_dat_data_d_2_72 = _RAND_200[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  in_rt_dat_data_d_2_73 = _RAND_201[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  in_rt_dat_data_d_2_74 = _RAND_202[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  in_rt_dat_data_d_2_75 = _RAND_203[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  in_rt_dat_data_d_2_76 = _RAND_204[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  in_rt_dat_data_d_2_77 = _RAND_205[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  in_rt_dat_data_d_2_78 = _RAND_206[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  in_rt_dat_data_d_2_79 = _RAND_207[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  in_rt_dat_data_d_2_80 = _RAND_208[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  in_rt_dat_data_d_2_81 = _RAND_209[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  in_rt_dat_data_d_2_82 = _RAND_210[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  in_rt_dat_data_d_2_83 = _RAND_211[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  in_rt_dat_data_d_2_84 = _RAND_212[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  in_rt_dat_data_d_2_85 = _RAND_213[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  in_rt_dat_data_d_2_86 = _RAND_214[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  in_rt_dat_data_d_2_87 = _RAND_215[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  in_rt_dat_data_d_2_88 = _RAND_216[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  in_rt_dat_data_d_2_89 = _RAND_217[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  in_rt_dat_data_d_2_90 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  in_rt_dat_data_d_2_91 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  in_rt_dat_data_d_2_92 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  in_rt_dat_data_d_2_93 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  in_rt_dat_data_d_2_94 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  in_rt_dat_data_d_2_95 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  in_rt_dat_data_d_2_96 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  in_rt_dat_data_d_2_97 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  in_rt_dat_data_d_2_98 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  in_rt_dat_data_d_2_99 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  in_rt_dat_data_d_2_100 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  in_rt_dat_data_d_2_101 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  in_rt_dat_data_d_2_102 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  in_rt_dat_data_d_2_103 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  in_rt_dat_data_d_2_104 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  in_rt_dat_data_d_2_105 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  in_rt_dat_data_d_2_106 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  in_rt_dat_data_d_2_107 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  in_rt_dat_data_d_2_108 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  in_rt_dat_data_d_2_109 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  in_rt_dat_data_d_2_110 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  in_rt_dat_data_d_2_111 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  in_rt_dat_data_d_2_112 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  in_rt_dat_data_d_2_113 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  in_rt_dat_data_d_2_114 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  in_rt_dat_data_d_2_115 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  in_rt_dat_data_d_2_116 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  in_rt_dat_data_d_2_117 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  in_rt_dat_data_d_2_118 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  in_rt_dat_data_d_2_119 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  in_rt_dat_data_d_2_120 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  in_rt_dat_data_d_2_121 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  in_rt_dat_data_d_2_122 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  in_rt_dat_data_d_2_123 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  in_rt_dat_data_d_2_124 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  in_rt_dat_data_d_2_125 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  in_rt_dat_data_d_2_126 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  in_rt_dat_data_d_2_127 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_0 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_1 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_2 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_3 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_4 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_5 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_6 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_7 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_8 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_9 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_10 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_11 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_12 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_13 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_14 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_15 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_16 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_17 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_18 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_19 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_20 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_21 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_22 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_23 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_24 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_25 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_26 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_27 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_28 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_29 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_30 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_31 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_32 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_33 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_34 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_35 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_36 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_37 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_38 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_39 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_40 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_41 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_42 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_43 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_44 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_45 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_46 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_47 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_48 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_49 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_50 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_51 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_52 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_53 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_54 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_55 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_56 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_57 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_58 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_59 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_60 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_61 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_62 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_63 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_64 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_65 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_66 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_67 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_68 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_69 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_70 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_71 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_72 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_73 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_74 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_75 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_76 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_77 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_78 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_79 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_80 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_81 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_82 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_83 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_84 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_85 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_86 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_87 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_88 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_89 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_90 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_91 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_92 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_93 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_94 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_95 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_96 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_97 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_98 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_99 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_100 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_101 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_102 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_103 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_104 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_105 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_106 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_107 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_108 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_109 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_110 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_111 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_112 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_113 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_114 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_115 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_116 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_117 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_118 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_119 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_120 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_121 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_122 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_123 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_124 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_125 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_126 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  in_rt_dat_mask_d_1_127 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_0 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_1 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_2 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_3 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_4 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_5 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_6 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_7 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_8 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_9 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_10 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_11 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_12 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_13 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_14 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_15 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_16 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_17 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_18 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_19 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_20 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_21 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_22 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_23 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_24 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_25 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_26 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_27 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_28 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_29 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_30 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_31 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_32 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_33 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_34 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_35 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_36 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_37 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_38 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_39 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_40 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_41 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_42 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_43 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_44 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_45 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_46 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_47 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_48 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_49 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_50 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_51 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_52 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_53 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_54 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_55 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_56 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_57 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_58 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_59 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_60 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_61 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_62 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_63 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_64 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_65 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_66 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_67 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_68 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_69 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_70 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_71 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_72 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_73 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_74 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_75 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_76 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_77 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_78 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_79 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_80 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_81 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_82 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_83 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_84 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_85 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_86 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_87 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_88 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_89 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_90 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_91 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_92 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_93 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_94 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_95 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_96 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_97 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_98 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_99 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_100 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_101 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_102 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_103 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_104 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_105 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_106 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_107 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_108 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_109 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_110 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_111 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_112 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_113 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_114 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_115 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_116 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_117 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_118 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_119 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_120 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_121 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_122 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_123 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_124 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_125 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_126 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  in_rt_dat_mask_d_2_127 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  in_rt_dat_pvld_d_1 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  in_rt_dat_pvld_d_2 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  in_rt_dat_pd_d_1 = _RAND_514[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  in_rt_dat_pd_d_2 = _RAND_515[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  in_rt_wt_data_d_1_0 = _RAND_516[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  in_rt_wt_data_d_1_1 = _RAND_517[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  in_rt_wt_data_d_1_2 = _RAND_518[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  in_rt_wt_data_d_1_3 = _RAND_519[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  in_rt_wt_data_d_1_4 = _RAND_520[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  in_rt_wt_data_d_1_5 = _RAND_521[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  in_rt_wt_data_d_1_6 = _RAND_522[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  in_rt_wt_data_d_1_7 = _RAND_523[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  in_rt_wt_data_d_1_8 = _RAND_524[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  in_rt_wt_data_d_1_9 = _RAND_525[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  in_rt_wt_data_d_1_10 = _RAND_526[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  in_rt_wt_data_d_1_11 = _RAND_527[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  in_rt_wt_data_d_1_12 = _RAND_528[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  in_rt_wt_data_d_1_13 = _RAND_529[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  in_rt_wt_data_d_1_14 = _RAND_530[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  in_rt_wt_data_d_1_15 = _RAND_531[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  in_rt_wt_data_d_1_16 = _RAND_532[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  in_rt_wt_data_d_1_17 = _RAND_533[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  in_rt_wt_data_d_1_18 = _RAND_534[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  in_rt_wt_data_d_1_19 = _RAND_535[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  in_rt_wt_data_d_1_20 = _RAND_536[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  in_rt_wt_data_d_1_21 = _RAND_537[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  in_rt_wt_data_d_1_22 = _RAND_538[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  in_rt_wt_data_d_1_23 = _RAND_539[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  in_rt_wt_data_d_1_24 = _RAND_540[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  in_rt_wt_data_d_1_25 = _RAND_541[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  in_rt_wt_data_d_1_26 = _RAND_542[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  in_rt_wt_data_d_1_27 = _RAND_543[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  in_rt_wt_data_d_1_28 = _RAND_544[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  in_rt_wt_data_d_1_29 = _RAND_545[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  in_rt_wt_data_d_1_30 = _RAND_546[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  in_rt_wt_data_d_1_31 = _RAND_547[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  in_rt_wt_data_d_1_32 = _RAND_548[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  in_rt_wt_data_d_1_33 = _RAND_549[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  in_rt_wt_data_d_1_34 = _RAND_550[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  in_rt_wt_data_d_1_35 = _RAND_551[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  in_rt_wt_data_d_1_36 = _RAND_552[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  in_rt_wt_data_d_1_37 = _RAND_553[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  in_rt_wt_data_d_1_38 = _RAND_554[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  in_rt_wt_data_d_1_39 = _RAND_555[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  in_rt_wt_data_d_1_40 = _RAND_556[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  in_rt_wt_data_d_1_41 = _RAND_557[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  in_rt_wt_data_d_1_42 = _RAND_558[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  in_rt_wt_data_d_1_43 = _RAND_559[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  in_rt_wt_data_d_1_44 = _RAND_560[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  in_rt_wt_data_d_1_45 = _RAND_561[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  in_rt_wt_data_d_1_46 = _RAND_562[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  in_rt_wt_data_d_1_47 = _RAND_563[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  in_rt_wt_data_d_1_48 = _RAND_564[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  in_rt_wt_data_d_1_49 = _RAND_565[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  in_rt_wt_data_d_1_50 = _RAND_566[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  in_rt_wt_data_d_1_51 = _RAND_567[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  in_rt_wt_data_d_1_52 = _RAND_568[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  in_rt_wt_data_d_1_53 = _RAND_569[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  in_rt_wt_data_d_1_54 = _RAND_570[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  in_rt_wt_data_d_1_55 = _RAND_571[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  in_rt_wt_data_d_1_56 = _RAND_572[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  in_rt_wt_data_d_1_57 = _RAND_573[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  in_rt_wt_data_d_1_58 = _RAND_574[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  in_rt_wt_data_d_1_59 = _RAND_575[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  in_rt_wt_data_d_1_60 = _RAND_576[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  in_rt_wt_data_d_1_61 = _RAND_577[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  in_rt_wt_data_d_1_62 = _RAND_578[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  in_rt_wt_data_d_1_63 = _RAND_579[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  in_rt_wt_data_d_1_64 = _RAND_580[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  in_rt_wt_data_d_1_65 = _RAND_581[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  in_rt_wt_data_d_1_66 = _RAND_582[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  in_rt_wt_data_d_1_67 = _RAND_583[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  in_rt_wt_data_d_1_68 = _RAND_584[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  in_rt_wt_data_d_1_69 = _RAND_585[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  in_rt_wt_data_d_1_70 = _RAND_586[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  in_rt_wt_data_d_1_71 = _RAND_587[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  in_rt_wt_data_d_1_72 = _RAND_588[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  in_rt_wt_data_d_1_73 = _RAND_589[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  in_rt_wt_data_d_1_74 = _RAND_590[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  in_rt_wt_data_d_1_75 = _RAND_591[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  in_rt_wt_data_d_1_76 = _RAND_592[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  in_rt_wt_data_d_1_77 = _RAND_593[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  in_rt_wt_data_d_1_78 = _RAND_594[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  in_rt_wt_data_d_1_79 = _RAND_595[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  in_rt_wt_data_d_1_80 = _RAND_596[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  in_rt_wt_data_d_1_81 = _RAND_597[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  in_rt_wt_data_d_1_82 = _RAND_598[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  in_rt_wt_data_d_1_83 = _RAND_599[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  in_rt_wt_data_d_1_84 = _RAND_600[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  in_rt_wt_data_d_1_85 = _RAND_601[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  in_rt_wt_data_d_1_86 = _RAND_602[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  in_rt_wt_data_d_1_87 = _RAND_603[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  in_rt_wt_data_d_1_88 = _RAND_604[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  in_rt_wt_data_d_1_89 = _RAND_605[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  in_rt_wt_data_d_1_90 = _RAND_606[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  in_rt_wt_data_d_1_91 = _RAND_607[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  in_rt_wt_data_d_1_92 = _RAND_608[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  in_rt_wt_data_d_1_93 = _RAND_609[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  in_rt_wt_data_d_1_94 = _RAND_610[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  in_rt_wt_data_d_1_95 = _RAND_611[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  in_rt_wt_data_d_1_96 = _RAND_612[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  in_rt_wt_data_d_1_97 = _RAND_613[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  in_rt_wt_data_d_1_98 = _RAND_614[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  in_rt_wt_data_d_1_99 = _RAND_615[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  in_rt_wt_data_d_1_100 = _RAND_616[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  in_rt_wt_data_d_1_101 = _RAND_617[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  in_rt_wt_data_d_1_102 = _RAND_618[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  in_rt_wt_data_d_1_103 = _RAND_619[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  in_rt_wt_data_d_1_104 = _RAND_620[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  in_rt_wt_data_d_1_105 = _RAND_621[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  in_rt_wt_data_d_1_106 = _RAND_622[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  in_rt_wt_data_d_1_107 = _RAND_623[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  in_rt_wt_data_d_1_108 = _RAND_624[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  in_rt_wt_data_d_1_109 = _RAND_625[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  in_rt_wt_data_d_1_110 = _RAND_626[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  in_rt_wt_data_d_1_111 = _RAND_627[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  in_rt_wt_data_d_1_112 = _RAND_628[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  in_rt_wt_data_d_1_113 = _RAND_629[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  in_rt_wt_data_d_1_114 = _RAND_630[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  in_rt_wt_data_d_1_115 = _RAND_631[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  in_rt_wt_data_d_1_116 = _RAND_632[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  in_rt_wt_data_d_1_117 = _RAND_633[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  in_rt_wt_data_d_1_118 = _RAND_634[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  in_rt_wt_data_d_1_119 = _RAND_635[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  in_rt_wt_data_d_1_120 = _RAND_636[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  in_rt_wt_data_d_1_121 = _RAND_637[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  in_rt_wt_data_d_1_122 = _RAND_638[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  in_rt_wt_data_d_1_123 = _RAND_639[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  in_rt_wt_data_d_1_124 = _RAND_640[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  in_rt_wt_data_d_1_125 = _RAND_641[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  in_rt_wt_data_d_1_126 = _RAND_642[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  in_rt_wt_data_d_1_127 = _RAND_643[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  in_rt_wt_data_d_2_0 = _RAND_644[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  in_rt_wt_data_d_2_1 = _RAND_645[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  in_rt_wt_data_d_2_2 = _RAND_646[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  in_rt_wt_data_d_2_3 = _RAND_647[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  in_rt_wt_data_d_2_4 = _RAND_648[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  in_rt_wt_data_d_2_5 = _RAND_649[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  in_rt_wt_data_d_2_6 = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  in_rt_wt_data_d_2_7 = _RAND_651[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  in_rt_wt_data_d_2_8 = _RAND_652[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  in_rt_wt_data_d_2_9 = _RAND_653[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  in_rt_wt_data_d_2_10 = _RAND_654[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  in_rt_wt_data_d_2_11 = _RAND_655[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  in_rt_wt_data_d_2_12 = _RAND_656[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  in_rt_wt_data_d_2_13 = _RAND_657[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  in_rt_wt_data_d_2_14 = _RAND_658[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  in_rt_wt_data_d_2_15 = _RAND_659[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  in_rt_wt_data_d_2_16 = _RAND_660[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  in_rt_wt_data_d_2_17 = _RAND_661[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  in_rt_wt_data_d_2_18 = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  in_rt_wt_data_d_2_19 = _RAND_663[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  in_rt_wt_data_d_2_20 = _RAND_664[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  in_rt_wt_data_d_2_21 = _RAND_665[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  in_rt_wt_data_d_2_22 = _RAND_666[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  in_rt_wt_data_d_2_23 = _RAND_667[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  in_rt_wt_data_d_2_24 = _RAND_668[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  in_rt_wt_data_d_2_25 = _RAND_669[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  in_rt_wt_data_d_2_26 = _RAND_670[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  in_rt_wt_data_d_2_27 = _RAND_671[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  in_rt_wt_data_d_2_28 = _RAND_672[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  in_rt_wt_data_d_2_29 = _RAND_673[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  in_rt_wt_data_d_2_30 = _RAND_674[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  in_rt_wt_data_d_2_31 = _RAND_675[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  in_rt_wt_data_d_2_32 = _RAND_676[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  in_rt_wt_data_d_2_33 = _RAND_677[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  in_rt_wt_data_d_2_34 = _RAND_678[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  in_rt_wt_data_d_2_35 = _RAND_679[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  in_rt_wt_data_d_2_36 = _RAND_680[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  in_rt_wt_data_d_2_37 = _RAND_681[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  in_rt_wt_data_d_2_38 = _RAND_682[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  in_rt_wt_data_d_2_39 = _RAND_683[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  in_rt_wt_data_d_2_40 = _RAND_684[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  in_rt_wt_data_d_2_41 = _RAND_685[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  in_rt_wt_data_d_2_42 = _RAND_686[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  in_rt_wt_data_d_2_43 = _RAND_687[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  in_rt_wt_data_d_2_44 = _RAND_688[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  in_rt_wt_data_d_2_45 = _RAND_689[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  in_rt_wt_data_d_2_46 = _RAND_690[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  in_rt_wt_data_d_2_47 = _RAND_691[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  in_rt_wt_data_d_2_48 = _RAND_692[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  in_rt_wt_data_d_2_49 = _RAND_693[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  in_rt_wt_data_d_2_50 = _RAND_694[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  in_rt_wt_data_d_2_51 = _RAND_695[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  in_rt_wt_data_d_2_52 = _RAND_696[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  in_rt_wt_data_d_2_53 = _RAND_697[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  in_rt_wt_data_d_2_54 = _RAND_698[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  in_rt_wt_data_d_2_55 = _RAND_699[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  in_rt_wt_data_d_2_56 = _RAND_700[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  in_rt_wt_data_d_2_57 = _RAND_701[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  in_rt_wt_data_d_2_58 = _RAND_702[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  in_rt_wt_data_d_2_59 = _RAND_703[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  in_rt_wt_data_d_2_60 = _RAND_704[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  in_rt_wt_data_d_2_61 = _RAND_705[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  in_rt_wt_data_d_2_62 = _RAND_706[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  in_rt_wt_data_d_2_63 = _RAND_707[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  in_rt_wt_data_d_2_64 = _RAND_708[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  in_rt_wt_data_d_2_65 = _RAND_709[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  in_rt_wt_data_d_2_66 = _RAND_710[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  in_rt_wt_data_d_2_67 = _RAND_711[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  in_rt_wt_data_d_2_68 = _RAND_712[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  in_rt_wt_data_d_2_69 = _RAND_713[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  in_rt_wt_data_d_2_70 = _RAND_714[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  in_rt_wt_data_d_2_71 = _RAND_715[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  in_rt_wt_data_d_2_72 = _RAND_716[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  in_rt_wt_data_d_2_73 = _RAND_717[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  in_rt_wt_data_d_2_74 = _RAND_718[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  in_rt_wt_data_d_2_75 = _RAND_719[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  in_rt_wt_data_d_2_76 = _RAND_720[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  in_rt_wt_data_d_2_77 = _RAND_721[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  in_rt_wt_data_d_2_78 = _RAND_722[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  in_rt_wt_data_d_2_79 = _RAND_723[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  in_rt_wt_data_d_2_80 = _RAND_724[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  in_rt_wt_data_d_2_81 = _RAND_725[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  in_rt_wt_data_d_2_82 = _RAND_726[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  in_rt_wt_data_d_2_83 = _RAND_727[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  in_rt_wt_data_d_2_84 = _RAND_728[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  in_rt_wt_data_d_2_85 = _RAND_729[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  in_rt_wt_data_d_2_86 = _RAND_730[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  in_rt_wt_data_d_2_87 = _RAND_731[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  in_rt_wt_data_d_2_88 = _RAND_732[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  in_rt_wt_data_d_2_89 = _RAND_733[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  in_rt_wt_data_d_2_90 = _RAND_734[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  in_rt_wt_data_d_2_91 = _RAND_735[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  in_rt_wt_data_d_2_92 = _RAND_736[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  in_rt_wt_data_d_2_93 = _RAND_737[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  in_rt_wt_data_d_2_94 = _RAND_738[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  in_rt_wt_data_d_2_95 = _RAND_739[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  in_rt_wt_data_d_2_96 = _RAND_740[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  in_rt_wt_data_d_2_97 = _RAND_741[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  in_rt_wt_data_d_2_98 = _RAND_742[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  in_rt_wt_data_d_2_99 = _RAND_743[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  in_rt_wt_data_d_2_100 = _RAND_744[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  in_rt_wt_data_d_2_101 = _RAND_745[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  in_rt_wt_data_d_2_102 = _RAND_746[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  in_rt_wt_data_d_2_103 = _RAND_747[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  in_rt_wt_data_d_2_104 = _RAND_748[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  in_rt_wt_data_d_2_105 = _RAND_749[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  in_rt_wt_data_d_2_106 = _RAND_750[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  in_rt_wt_data_d_2_107 = _RAND_751[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  in_rt_wt_data_d_2_108 = _RAND_752[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  in_rt_wt_data_d_2_109 = _RAND_753[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  in_rt_wt_data_d_2_110 = _RAND_754[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  in_rt_wt_data_d_2_111 = _RAND_755[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  in_rt_wt_data_d_2_112 = _RAND_756[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  in_rt_wt_data_d_2_113 = _RAND_757[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  in_rt_wt_data_d_2_114 = _RAND_758[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  in_rt_wt_data_d_2_115 = _RAND_759[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  in_rt_wt_data_d_2_116 = _RAND_760[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  in_rt_wt_data_d_2_117 = _RAND_761[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  in_rt_wt_data_d_2_118 = _RAND_762[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  in_rt_wt_data_d_2_119 = _RAND_763[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  in_rt_wt_data_d_2_120 = _RAND_764[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  in_rt_wt_data_d_2_121 = _RAND_765[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  in_rt_wt_data_d_2_122 = _RAND_766[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  in_rt_wt_data_d_2_123 = _RAND_767[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  in_rt_wt_data_d_2_124 = _RAND_768[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  in_rt_wt_data_d_2_125 = _RAND_769[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  in_rt_wt_data_d_2_126 = _RAND_770[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  in_rt_wt_data_d_2_127 = _RAND_771[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_0 = _RAND_772[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_1 = _RAND_773[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_2 = _RAND_774[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_3 = _RAND_775[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_4 = _RAND_776[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_5 = _RAND_777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_6 = _RAND_778[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_7 = _RAND_779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_8 = _RAND_780[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_9 = _RAND_781[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_10 = _RAND_782[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_11 = _RAND_783[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_12 = _RAND_784[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_13 = _RAND_785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_14 = _RAND_786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_15 = _RAND_787[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_16 = _RAND_788[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_17 = _RAND_789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_18 = _RAND_790[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_19 = _RAND_791[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_20 = _RAND_792[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_21 = _RAND_793[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_22 = _RAND_794[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_23 = _RAND_795[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_24 = _RAND_796[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_25 = _RAND_797[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_26 = _RAND_798[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_27 = _RAND_799[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_28 = _RAND_800[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_29 = _RAND_801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_30 = _RAND_802[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_31 = _RAND_803[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_32 = _RAND_804[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_33 = _RAND_805[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_34 = _RAND_806[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_35 = _RAND_807[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_36 = _RAND_808[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_37 = _RAND_809[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_38 = _RAND_810[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_39 = _RAND_811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_40 = _RAND_812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_41 = _RAND_813[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_42 = _RAND_814[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_43 = _RAND_815[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_44 = _RAND_816[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_45 = _RAND_817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_46 = _RAND_818[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_47 = _RAND_819[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_48 = _RAND_820[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_49 = _RAND_821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_50 = _RAND_822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_51 = _RAND_823[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_52 = _RAND_824[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_53 = _RAND_825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_54 = _RAND_826[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_55 = _RAND_827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_56 = _RAND_828[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_57 = _RAND_829[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_58 = _RAND_830[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_59 = _RAND_831[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_60 = _RAND_832[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_61 = _RAND_833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_62 = _RAND_834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_63 = _RAND_835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_64 = _RAND_836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_65 = _RAND_837[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_66 = _RAND_838[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_67 = _RAND_839[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_68 = _RAND_840[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_69 = _RAND_841[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_70 = _RAND_842[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_71 = _RAND_843[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_72 = _RAND_844[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_73 = _RAND_845[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_74 = _RAND_846[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_75 = _RAND_847[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_76 = _RAND_848[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_77 = _RAND_849[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_78 = _RAND_850[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_79 = _RAND_851[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_80 = _RAND_852[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_81 = _RAND_853[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_82 = _RAND_854[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_83 = _RAND_855[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_84 = _RAND_856[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_85 = _RAND_857[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_86 = _RAND_858[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_87 = _RAND_859[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_88 = _RAND_860[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_89 = _RAND_861[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_90 = _RAND_862[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_91 = _RAND_863[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_92 = _RAND_864[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_93 = _RAND_865[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_94 = _RAND_866[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_95 = _RAND_867[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_96 = _RAND_868[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_97 = _RAND_869[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_98 = _RAND_870[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_99 = _RAND_871[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_100 = _RAND_872[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_101 = _RAND_873[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_102 = _RAND_874[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_103 = _RAND_875[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_104 = _RAND_876[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_105 = _RAND_877[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_106 = _RAND_878[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_107 = _RAND_879[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_108 = _RAND_880[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_109 = _RAND_881[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_110 = _RAND_882[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_111 = _RAND_883[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_112 = _RAND_884[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_113 = _RAND_885[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_114 = _RAND_886[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_115 = _RAND_887[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_116 = _RAND_888[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_117 = _RAND_889[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_118 = _RAND_890[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_119 = _RAND_891[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_120 = _RAND_892[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_121 = _RAND_893[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_122 = _RAND_894[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_123 = _RAND_895[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_124 = _RAND_896[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_125 = _RAND_897[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_126 = _RAND_898[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  in_rt_wt_mask_d_1_127 = _RAND_899[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_0 = _RAND_900[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_1 = _RAND_901[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_2 = _RAND_902[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_3 = _RAND_903[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_4 = _RAND_904[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_5 = _RAND_905[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_6 = _RAND_906[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_7 = _RAND_907[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_8 = _RAND_908[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_9 = _RAND_909[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_10 = _RAND_910[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_11 = _RAND_911[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_12 = _RAND_912[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_13 = _RAND_913[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_14 = _RAND_914[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_15 = _RAND_915[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_16 = _RAND_916[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_17 = _RAND_917[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_18 = _RAND_918[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_19 = _RAND_919[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_20 = _RAND_920[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_21 = _RAND_921[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_22 = _RAND_922[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_23 = _RAND_923[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_24 = _RAND_924[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_25 = _RAND_925[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_26 = _RAND_926[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_27 = _RAND_927[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_28 = _RAND_928[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_29 = _RAND_929[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_30 = _RAND_930[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_31 = _RAND_931[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_32 = _RAND_932[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_33 = _RAND_933[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_34 = _RAND_934[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_35 = _RAND_935[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_36 = _RAND_936[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_37 = _RAND_937[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_38 = _RAND_938[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_39 = _RAND_939[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_40 = _RAND_940[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_41 = _RAND_941[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_42 = _RAND_942[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_43 = _RAND_943[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_44 = _RAND_944[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_45 = _RAND_945[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_46 = _RAND_946[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_47 = _RAND_947[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_48 = _RAND_948[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_49 = _RAND_949[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_50 = _RAND_950[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_51 = _RAND_951[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_52 = _RAND_952[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_53 = _RAND_953[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_54 = _RAND_954[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_55 = _RAND_955[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_56 = _RAND_956[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_57 = _RAND_957[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_58 = _RAND_958[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_59 = _RAND_959[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_60 = _RAND_960[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_61 = _RAND_961[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_62 = _RAND_962[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_63 = _RAND_963[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_64 = _RAND_964[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_65 = _RAND_965[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_66 = _RAND_966[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_67 = _RAND_967[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_68 = _RAND_968[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_69 = _RAND_969[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_70 = _RAND_970[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_71 = _RAND_971[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_72 = _RAND_972[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_73 = _RAND_973[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_74 = _RAND_974[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_75 = _RAND_975[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_76 = _RAND_976[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_77 = _RAND_977[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_78 = _RAND_978[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_79 = _RAND_979[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_80 = _RAND_980[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_81 = _RAND_981[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_82 = _RAND_982[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_83 = _RAND_983[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_84 = _RAND_984[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_85 = _RAND_985[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_86 = _RAND_986[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_87 = _RAND_987[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_88 = _RAND_988[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_89 = _RAND_989[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_90 = _RAND_990[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_91 = _RAND_991[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_92 = _RAND_992[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_93 = _RAND_993[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_94 = _RAND_994[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_95 = _RAND_995[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_96 = _RAND_996[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_97 = _RAND_997[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_98 = _RAND_998[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_99 = _RAND_999[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_100 = _RAND_1000[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_101 = _RAND_1001[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_102 = _RAND_1002[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_103 = _RAND_1003[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_104 = _RAND_1004[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_105 = _RAND_1005[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_106 = _RAND_1006[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_107 = _RAND_1007[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_108 = _RAND_1008[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_109 = _RAND_1009[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_110 = _RAND_1010[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_111 = _RAND_1011[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_112 = _RAND_1012[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_113 = _RAND_1013[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_114 = _RAND_1014[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_115 = _RAND_1015[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_116 = _RAND_1016[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_117 = _RAND_1017[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_118 = _RAND_1018[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_119 = _RAND_1019[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_120 = _RAND_1020[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_121 = _RAND_1021[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_122 = _RAND_1022[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_123 = _RAND_1023[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_124 = _RAND_1024[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_125 = _RAND_1025[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_126 = _RAND_1026[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  in_rt_wt_mask_d_2_127 = _RAND_1027[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  in_rt_wt_pvld_d_1 = _RAND_1028[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  in_rt_wt_pvld_d_2 = _RAND_1029[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  in_rt_wt_sel_d_1_0 = _RAND_1030[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  in_rt_wt_sel_d_2_0 = _RAND_1031[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_sc2mac_dat_mask_0) begin
      in_rt_dat_data_d_1_0 <= io_sc2mac_dat_data_0;
    end
    if (io_sc2mac_dat_mask_1) begin
      in_rt_dat_data_d_1_1 <= io_sc2mac_dat_data_1;
    end
    if (io_sc2mac_dat_mask_2) begin
      in_rt_dat_data_d_1_2 <= io_sc2mac_dat_data_2;
    end
    if (io_sc2mac_dat_mask_3) begin
      in_rt_dat_data_d_1_3 <= io_sc2mac_dat_data_3;
    end
    if (io_sc2mac_dat_mask_4) begin
      in_rt_dat_data_d_1_4 <= io_sc2mac_dat_data_4;
    end
    if (io_sc2mac_dat_mask_5) begin
      in_rt_dat_data_d_1_5 <= io_sc2mac_dat_data_5;
    end
    if (io_sc2mac_dat_mask_6) begin
      in_rt_dat_data_d_1_6 <= io_sc2mac_dat_data_6;
    end
    if (io_sc2mac_dat_mask_7) begin
      in_rt_dat_data_d_1_7 <= io_sc2mac_dat_data_7;
    end
    if (io_sc2mac_dat_mask_8) begin
      in_rt_dat_data_d_1_8 <= io_sc2mac_dat_data_8;
    end
    if (io_sc2mac_dat_mask_9) begin
      in_rt_dat_data_d_1_9 <= io_sc2mac_dat_data_9;
    end
    if (io_sc2mac_dat_mask_10) begin
      in_rt_dat_data_d_1_10 <= io_sc2mac_dat_data_10;
    end
    if (io_sc2mac_dat_mask_11) begin
      in_rt_dat_data_d_1_11 <= io_sc2mac_dat_data_11;
    end
    if (io_sc2mac_dat_mask_12) begin
      in_rt_dat_data_d_1_12 <= io_sc2mac_dat_data_12;
    end
    if (io_sc2mac_dat_mask_13) begin
      in_rt_dat_data_d_1_13 <= io_sc2mac_dat_data_13;
    end
    if (io_sc2mac_dat_mask_14) begin
      in_rt_dat_data_d_1_14 <= io_sc2mac_dat_data_14;
    end
    if (io_sc2mac_dat_mask_15) begin
      in_rt_dat_data_d_1_15 <= io_sc2mac_dat_data_15;
    end
    if (io_sc2mac_dat_mask_16) begin
      in_rt_dat_data_d_1_16 <= io_sc2mac_dat_data_16;
    end
    if (io_sc2mac_dat_mask_17) begin
      in_rt_dat_data_d_1_17 <= io_sc2mac_dat_data_17;
    end
    if (io_sc2mac_dat_mask_18) begin
      in_rt_dat_data_d_1_18 <= io_sc2mac_dat_data_18;
    end
    if (io_sc2mac_dat_mask_19) begin
      in_rt_dat_data_d_1_19 <= io_sc2mac_dat_data_19;
    end
    if (io_sc2mac_dat_mask_20) begin
      in_rt_dat_data_d_1_20 <= io_sc2mac_dat_data_20;
    end
    if (io_sc2mac_dat_mask_21) begin
      in_rt_dat_data_d_1_21 <= io_sc2mac_dat_data_21;
    end
    if (io_sc2mac_dat_mask_22) begin
      in_rt_dat_data_d_1_22 <= io_sc2mac_dat_data_22;
    end
    if (io_sc2mac_dat_mask_23) begin
      in_rt_dat_data_d_1_23 <= io_sc2mac_dat_data_23;
    end
    if (io_sc2mac_dat_mask_24) begin
      in_rt_dat_data_d_1_24 <= io_sc2mac_dat_data_24;
    end
    if (io_sc2mac_dat_mask_25) begin
      in_rt_dat_data_d_1_25 <= io_sc2mac_dat_data_25;
    end
    if (io_sc2mac_dat_mask_26) begin
      in_rt_dat_data_d_1_26 <= io_sc2mac_dat_data_26;
    end
    if (io_sc2mac_dat_mask_27) begin
      in_rt_dat_data_d_1_27 <= io_sc2mac_dat_data_27;
    end
    if (io_sc2mac_dat_mask_28) begin
      in_rt_dat_data_d_1_28 <= io_sc2mac_dat_data_28;
    end
    if (io_sc2mac_dat_mask_29) begin
      in_rt_dat_data_d_1_29 <= io_sc2mac_dat_data_29;
    end
    if (io_sc2mac_dat_mask_30) begin
      in_rt_dat_data_d_1_30 <= io_sc2mac_dat_data_30;
    end
    if (io_sc2mac_dat_mask_31) begin
      in_rt_dat_data_d_1_31 <= io_sc2mac_dat_data_31;
    end
    if (io_sc2mac_dat_mask_32) begin
      in_rt_dat_data_d_1_32 <= io_sc2mac_dat_data_32;
    end
    if (io_sc2mac_dat_mask_33) begin
      in_rt_dat_data_d_1_33 <= io_sc2mac_dat_data_33;
    end
    if (io_sc2mac_dat_mask_34) begin
      in_rt_dat_data_d_1_34 <= io_sc2mac_dat_data_34;
    end
    if (io_sc2mac_dat_mask_35) begin
      in_rt_dat_data_d_1_35 <= io_sc2mac_dat_data_35;
    end
    if (io_sc2mac_dat_mask_36) begin
      in_rt_dat_data_d_1_36 <= io_sc2mac_dat_data_36;
    end
    if (io_sc2mac_dat_mask_37) begin
      in_rt_dat_data_d_1_37 <= io_sc2mac_dat_data_37;
    end
    if (io_sc2mac_dat_mask_38) begin
      in_rt_dat_data_d_1_38 <= io_sc2mac_dat_data_38;
    end
    if (io_sc2mac_dat_mask_39) begin
      in_rt_dat_data_d_1_39 <= io_sc2mac_dat_data_39;
    end
    if (io_sc2mac_dat_mask_40) begin
      in_rt_dat_data_d_1_40 <= io_sc2mac_dat_data_40;
    end
    if (io_sc2mac_dat_mask_41) begin
      in_rt_dat_data_d_1_41 <= io_sc2mac_dat_data_41;
    end
    if (io_sc2mac_dat_mask_42) begin
      in_rt_dat_data_d_1_42 <= io_sc2mac_dat_data_42;
    end
    if (io_sc2mac_dat_mask_43) begin
      in_rt_dat_data_d_1_43 <= io_sc2mac_dat_data_43;
    end
    if (io_sc2mac_dat_mask_44) begin
      in_rt_dat_data_d_1_44 <= io_sc2mac_dat_data_44;
    end
    if (io_sc2mac_dat_mask_45) begin
      in_rt_dat_data_d_1_45 <= io_sc2mac_dat_data_45;
    end
    if (io_sc2mac_dat_mask_46) begin
      in_rt_dat_data_d_1_46 <= io_sc2mac_dat_data_46;
    end
    if (io_sc2mac_dat_mask_47) begin
      in_rt_dat_data_d_1_47 <= io_sc2mac_dat_data_47;
    end
    if (io_sc2mac_dat_mask_48) begin
      in_rt_dat_data_d_1_48 <= io_sc2mac_dat_data_48;
    end
    if (io_sc2mac_dat_mask_49) begin
      in_rt_dat_data_d_1_49 <= io_sc2mac_dat_data_49;
    end
    if (io_sc2mac_dat_mask_50) begin
      in_rt_dat_data_d_1_50 <= io_sc2mac_dat_data_50;
    end
    if (io_sc2mac_dat_mask_51) begin
      in_rt_dat_data_d_1_51 <= io_sc2mac_dat_data_51;
    end
    if (io_sc2mac_dat_mask_52) begin
      in_rt_dat_data_d_1_52 <= io_sc2mac_dat_data_52;
    end
    if (io_sc2mac_dat_mask_53) begin
      in_rt_dat_data_d_1_53 <= io_sc2mac_dat_data_53;
    end
    if (io_sc2mac_dat_mask_54) begin
      in_rt_dat_data_d_1_54 <= io_sc2mac_dat_data_54;
    end
    if (io_sc2mac_dat_mask_55) begin
      in_rt_dat_data_d_1_55 <= io_sc2mac_dat_data_55;
    end
    if (io_sc2mac_dat_mask_56) begin
      in_rt_dat_data_d_1_56 <= io_sc2mac_dat_data_56;
    end
    if (io_sc2mac_dat_mask_57) begin
      in_rt_dat_data_d_1_57 <= io_sc2mac_dat_data_57;
    end
    if (io_sc2mac_dat_mask_58) begin
      in_rt_dat_data_d_1_58 <= io_sc2mac_dat_data_58;
    end
    if (io_sc2mac_dat_mask_59) begin
      in_rt_dat_data_d_1_59 <= io_sc2mac_dat_data_59;
    end
    if (io_sc2mac_dat_mask_60) begin
      in_rt_dat_data_d_1_60 <= io_sc2mac_dat_data_60;
    end
    if (io_sc2mac_dat_mask_61) begin
      in_rt_dat_data_d_1_61 <= io_sc2mac_dat_data_61;
    end
    if (io_sc2mac_dat_mask_62) begin
      in_rt_dat_data_d_1_62 <= io_sc2mac_dat_data_62;
    end
    if (io_sc2mac_dat_mask_63) begin
      in_rt_dat_data_d_1_63 <= io_sc2mac_dat_data_63;
    end
    if (io_sc2mac_dat_mask_64) begin
      in_rt_dat_data_d_1_64 <= io_sc2mac_dat_data_64;
    end
    if (io_sc2mac_dat_mask_65) begin
      in_rt_dat_data_d_1_65 <= io_sc2mac_dat_data_65;
    end
    if (io_sc2mac_dat_mask_66) begin
      in_rt_dat_data_d_1_66 <= io_sc2mac_dat_data_66;
    end
    if (io_sc2mac_dat_mask_67) begin
      in_rt_dat_data_d_1_67 <= io_sc2mac_dat_data_67;
    end
    if (io_sc2mac_dat_mask_68) begin
      in_rt_dat_data_d_1_68 <= io_sc2mac_dat_data_68;
    end
    if (io_sc2mac_dat_mask_69) begin
      in_rt_dat_data_d_1_69 <= io_sc2mac_dat_data_69;
    end
    if (io_sc2mac_dat_mask_70) begin
      in_rt_dat_data_d_1_70 <= io_sc2mac_dat_data_70;
    end
    if (io_sc2mac_dat_mask_71) begin
      in_rt_dat_data_d_1_71 <= io_sc2mac_dat_data_71;
    end
    if (io_sc2mac_dat_mask_72) begin
      in_rt_dat_data_d_1_72 <= io_sc2mac_dat_data_72;
    end
    if (io_sc2mac_dat_mask_73) begin
      in_rt_dat_data_d_1_73 <= io_sc2mac_dat_data_73;
    end
    if (io_sc2mac_dat_mask_74) begin
      in_rt_dat_data_d_1_74 <= io_sc2mac_dat_data_74;
    end
    if (io_sc2mac_dat_mask_75) begin
      in_rt_dat_data_d_1_75 <= io_sc2mac_dat_data_75;
    end
    if (io_sc2mac_dat_mask_76) begin
      in_rt_dat_data_d_1_76 <= io_sc2mac_dat_data_76;
    end
    if (io_sc2mac_dat_mask_77) begin
      in_rt_dat_data_d_1_77 <= io_sc2mac_dat_data_77;
    end
    if (io_sc2mac_dat_mask_78) begin
      in_rt_dat_data_d_1_78 <= io_sc2mac_dat_data_78;
    end
    if (io_sc2mac_dat_mask_79) begin
      in_rt_dat_data_d_1_79 <= io_sc2mac_dat_data_79;
    end
    if (io_sc2mac_dat_mask_80) begin
      in_rt_dat_data_d_1_80 <= io_sc2mac_dat_data_80;
    end
    if (io_sc2mac_dat_mask_81) begin
      in_rt_dat_data_d_1_81 <= io_sc2mac_dat_data_81;
    end
    if (io_sc2mac_dat_mask_82) begin
      in_rt_dat_data_d_1_82 <= io_sc2mac_dat_data_82;
    end
    if (io_sc2mac_dat_mask_83) begin
      in_rt_dat_data_d_1_83 <= io_sc2mac_dat_data_83;
    end
    if (io_sc2mac_dat_mask_84) begin
      in_rt_dat_data_d_1_84 <= io_sc2mac_dat_data_84;
    end
    if (io_sc2mac_dat_mask_85) begin
      in_rt_dat_data_d_1_85 <= io_sc2mac_dat_data_85;
    end
    if (io_sc2mac_dat_mask_86) begin
      in_rt_dat_data_d_1_86 <= io_sc2mac_dat_data_86;
    end
    if (io_sc2mac_dat_mask_87) begin
      in_rt_dat_data_d_1_87 <= io_sc2mac_dat_data_87;
    end
    if (io_sc2mac_dat_mask_88) begin
      in_rt_dat_data_d_1_88 <= io_sc2mac_dat_data_88;
    end
    if (io_sc2mac_dat_mask_89) begin
      in_rt_dat_data_d_1_89 <= io_sc2mac_dat_data_89;
    end
    if (io_sc2mac_dat_mask_90) begin
      in_rt_dat_data_d_1_90 <= io_sc2mac_dat_data_90;
    end
    if (io_sc2mac_dat_mask_91) begin
      in_rt_dat_data_d_1_91 <= io_sc2mac_dat_data_91;
    end
    if (io_sc2mac_dat_mask_92) begin
      in_rt_dat_data_d_1_92 <= io_sc2mac_dat_data_92;
    end
    if (io_sc2mac_dat_mask_93) begin
      in_rt_dat_data_d_1_93 <= io_sc2mac_dat_data_93;
    end
    if (io_sc2mac_dat_mask_94) begin
      in_rt_dat_data_d_1_94 <= io_sc2mac_dat_data_94;
    end
    if (io_sc2mac_dat_mask_95) begin
      in_rt_dat_data_d_1_95 <= io_sc2mac_dat_data_95;
    end
    if (io_sc2mac_dat_mask_96) begin
      in_rt_dat_data_d_1_96 <= io_sc2mac_dat_data_96;
    end
    if (io_sc2mac_dat_mask_97) begin
      in_rt_dat_data_d_1_97 <= io_sc2mac_dat_data_97;
    end
    if (io_sc2mac_dat_mask_98) begin
      in_rt_dat_data_d_1_98 <= io_sc2mac_dat_data_98;
    end
    if (io_sc2mac_dat_mask_99) begin
      in_rt_dat_data_d_1_99 <= io_sc2mac_dat_data_99;
    end
    if (io_sc2mac_dat_mask_100) begin
      in_rt_dat_data_d_1_100 <= io_sc2mac_dat_data_100;
    end
    if (io_sc2mac_dat_mask_101) begin
      in_rt_dat_data_d_1_101 <= io_sc2mac_dat_data_101;
    end
    if (io_sc2mac_dat_mask_102) begin
      in_rt_dat_data_d_1_102 <= io_sc2mac_dat_data_102;
    end
    if (io_sc2mac_dat_mask_103) begin
      in_rt_dat_data_d_1_103 <= io_sc2mac_dat_data_103;
    end
    if (io_sc2mac_dat_mask_104) begin
      in_rt_dat_data_d_1_104 <= io_sc2mac_dat_data_104;
    end
    if (io_sc2mac_dat_mask_105) begin
      in_rt_dat_data_d_1_105 <= io_sc2mac_dat_data_105;
    end
    if (io_sc2mac_dat_mask_106) begin
      in_rt_dat_data_d_1_106 <= io_sc2mac_dat_data_106;
    end
    if (io_sc2mac_dat_mask_107) begin
      in_rt_dat_data_d_1_107 <= io_sc2mac_dat_data_107;
    end
    if (io_sc2mac_dat_mask_108) begin
      in_rt_dat_data_d_1_108 <= io_sc2mac_dat_data_108;
    end
    if (io_sc2mac_dat_mask_109) begin
      in_rt_dat_data_d_1_109 <= io_sc2mac_dat_data_109;
    end
    if (io_sc2mac_dat_mask_110) begin
      in_rt_dat_data_d_1_110 <= io_sc2mac_dat_data_110;
    end
    if (io_sc2mac_dat_mask_111) begin
      in_rt_dat_data_d_1_111 <= io_sc2mac_dat_data_111;
    end
    if (io_sc2mac_dat_mask_112) begin
      in_rt_dat_data_d_1_112 <= io_sc2mac_dat_data_112;
    end
    if (io_sc2mac_dat_mask_113) begin
      in_rt_dat_data_d_1_113 <= io_sc2mac_dat_data_113;
    end
    if (io_sc2mac_dat_mask_114) begin
      in_rt_dat_data_d_1_114 <= io_sc2mac_dat_data_114;
    end
    if (io_sc2mac_dat_mask_115) begin
      in_rt_dat_data_d_1_115 <= io_sc2mac_dat_data_115;
    end
    if (io_sc2mac_dat_mask_116) begin
      in_rt_dat_data_d_1_116 <= io_sc2mac_dat_data_116;
    end
    if (io_sc2mac_dat_mask_117) begin
      in_rt_dat_data_d_1_117 <= io_sc2mac_dat_data_117;
    end
    if (io_sc2mac_dat_mask_118) begin
      in_rt_dat_data_d_1_118 <= io_sc2mac_dat_data_118;
    end
    if (io_sc2mac_dat_mask_119) begin
      in_rt_dat_data_d_1_119 <= io_sc2mac_dat_data_119;
    end
    if (io_sc2mac_dat_mask_120) begin
      in_rt_dat_data_d_1_120 <= io_sc2mac_dat_data_120;
    end
    if (io_sc2mac_dat_mask_121) begin
      in_rt_dat_data_d_1_121 <= io_sc2mac_dat_data_121;
    end
    if (io_sc2mac_dat_mask_122) begin
      in_rt_dat_data_d_1_122 <= io_sc2mac_dat_data_122;
    end
    if (io_sc2mac_dat_mask_123) begin
      in_rt_dat_data_d_1_123 <= io_sc2mac_dat_data_123;
    end
    if (io_sc2mac_dat_mask_124) begin
      in_rt_dat_data_d_1_124 <= io_sc2mac_dat_data_124;
    end
    if (io_sc2mac_dat_mask_125) begin
      in_rt_dat_data_d_1_125 <= io_sc2mac_dat_data_125;
    end
    if (io_sc2mac_dat_mask_126) begin
      in_rt_dat_data_d_1_126 <= io_sc2mac_dat_data_126;
    end
    if (io_sc2mac_dat_mask_127) begin
      in_rt_dat_data_d_1_127 <= io_sc2mac_dat_data_127;
    end
    if (in_rt_dat_mask_d_1_0) begin
      in_rt_dat_data_d_2_0 <= in_rt_dat_data_d_1_0;
    end
    if (in_rt_dat_mask_d_1_1) begin
      in_rt_dat_data_d_2_1 <= in_rt_dat_data_d_1_1;
    end
    if (in_rt_dat_mask_d_1_2) begin
      in_rt_dat_data_d_2_2 <= in_rt_dat_data_d_1_2;
    end
    if (in_rt_dat_mask_d_1_3) begin
      in_rt_dat_data_d_2_3 <= in_rt_dat_data_d_1_3;
    end
    if (in_rt_dat_mask_d_1_4) begin
      in_rt_dat_data_d_2_4 <= in_rt_dat_data_d_1_4;
    end
    if (in_rt_dat_mask_d_1_5) begin
      in_rt_dat_data_d_2_5 <= in_rt_dat_data_d_1_5;
    end
    if (in_rt_dat_mask_d_1_6) begin
      in_rt_dat_data_d_2_6 <= in_rt_dat_data_d_1_6;
    end
    if (in_rt_dat_mask_d_1_7) begin
      in_rt_dat_data_d_2_7 <= in_rt_dat_data_d_1_7;
    end
    if (in_rt_dat_mask_d_1_8) begin
      in_rt_dat_data_d_2_8 <= in_rt_dat_data_d_1_8;
    end
    if (in_rt_dat_mask_d_1_9) begin
      in_rt_dat_data_d_2_9 <= in_rt_dat_data_d_1_9;
    end
    if (in_rt_dat_mask_d_1_10) begin
      in_rt_dat_data_d_2_10 <= in_rt_dat_data_d_1_10;
    end
    if (in_rt_dat_mask_d_1_11) begin
      in_rt_dat_data_d_2_11 <= in_rt_dat_data_d_1_11;
    end
    if (in_rt_dat_mask_d_1_12) begin
      in_rt_dat_data_d_2_12 <= in_rt_dat_data_d_1_12;
    end
    if (in_rt_dat_mask_d_1_13) begin
      in_rt_dat_data_d_2_13 <= in_rt_dat_data_d_1_13;
    end
    if (in_rt_dat_mask_d_1_14) begin
      in_rt_dat_data_d_2_14 <= in_rt_dat_data_d_1_14;
    end
    if (in_rt_dat_mask_d_1_15) begin
      in_rt_dat_data_d_2_15 <= in_rt_dat_data_d_1_15;
    end
    if (in_rt_dat_mask_d_1_16) begin
      in_rt_dat_data_d_2_16 <= in_rt_dat_data_d_1_16;
    end
    if (in_rt_dat_mask_d_1_17) begin
      in_rt_dat_data_d_2_17 <= in_rt_dat_data_d_1_17;
    end
    if (in_rt_dat_mask_d_1_18) begin
      in_rt_dat_data_d_2_18 <= in_rt_dat_data_d_1_18;
    end
    if (in_rt_dat_mask_d_1_19) begin
      in_rt_dat_data_d_2_19 <= in_rt_dat_data_d_1_19;
    end
    if (in_rt_dat_mask_d_1_20) begin
      in_rt_dat_data_d_2_20 <= in_rt_dat_data_d_1_20;
    end
    if (in_rt_dat_mask_d_1_21) begin
      in_rt_dat_data_d_2_21 <= in_rt_dat_data_d_1_21;
    end
    if (in_rt_dat_mask_d_1_22) begin
      in_rt_dat_data_d_2_22 <= in_rt_dat_data_d_1_22;
    end
    if (in_rt_dat_mask_d_1_23) begin
      in_rt_dat_data_d_2_23 <= in_rt_dat_data_d_1_23;
    end
    if (in_rt_dat_mask_d_1_24) begin
      in_rt_dat_data_d_2_24 <= in_rt_dat_data_d_1_24;
    end
    if (in_rt_dat_mask_d_1_25) begin
      in_rt_dat_data_d_2_25 <= in_rt_dat_data_d_1_25;
    end
    if (in_rt_dat_mask_d_1_26) begin
      in_rt_dat_data_d_2_26 <= in_rt_dat_data_d_1_26;
    end
    if (in_rt_dat_mask_d_1_27) begin
      in_rt_dat_data_d_2_27 <= in_rt_dat_data_d_1_27;
    end
    if (in_rt_dat_mask_d_1_28) begin
      in_rt_dat_data_d_2_28 <= in_rt_dat_data_d_1_28;
    end
    if (in_rt_dat_mask_d_1_29) begin
      in_rt_dat_data_d_2_29 <= in_rt_dat_data_d_1_29;
    end
    if (in_rt_dat_mask_d_1_30) begin
      in_rt_dat_data_d_2_30 <= in_rt_dat_data_d_1_30;
    end
    if (in_rt_dat_mask_d_1_31) begin
      in_rt_dat_data_d_2_31 <= in_rt_dat_data_d_1_31;
    end
    if (in_rt_dat_mask_d_1_32) begin
      in_rt_dat_data_d_2_32 <= in_rt_dat_data_d_1_32;
    end
    if (in_rt_dat_mask_d_1_33) begin
      in_rt_dat_data_d_2_33 <= in_rt_dat_data_d_1_33;
    end
    if (in_rt_dat_mask_d_1_34) begin
      in_rt_dat_data_d_2_34 <= in_rt_dat_data_d_1_34;
    end
    if (in_rt_dat_mask_d_1_35) begin
      in_rt_dat_data_d_2_35 <= in_rt_dat_data_d_1_35;
    end
    if (in_rt_dat_mask_d_1_36) begin
      in_rt_dat_data_d_2_36 <= in_rt_dat_data_d_1_36;
    end
    if (in_rt_dat_mask_d_1_37) begin
      in_rt_dat_data_d_2_37 <= in_rt_dat_data_d_1_37;
    end
    if (in_rt_dat_mask_d_1_38) begin
      in_rt_dat_data_d_2_38 <= in_rt_dat_data_d_1_38;
    end
    if (in_rt_dat_mask_d_1_39) begin
      in_rt_dat_data_d_2_39 <= in_rt_dat_data_d_1_39;
    end
    if (in_rt_dat_mask_d_1_40) begin
      in_rt_dat_data_d_2_40 <= in_rt_dat_data_d_1_40;
    end
    if (in_rt_dat_mask_d_1_41) begin
      in_rt_dat_data_d_2_41 <= in_rt_dat_data_d_1_41;
    end
    if (in_rt_dat_mask_d_1_42) begin
      in_rt_dat_data_d_2_42 <= in_rt_dat_data_d_1_42;
    end
    if (in_rt_dat_mask_d_1_43) begin
      in_rt_dat_data_d_2_43 <= in_rt_dat_data_d_1_43;
    end
    if (in_rt_dat_mask_d_1_44) begin
      in_rt_dat_data_d_2_44 <= in_rt_dat_data_d_1_44;
    end
    if (in_rt_dat_mask_d_1_45) begin
      in_rt_dat_data_d_2_45 <= in_rt_dat_data_d_1_45;
    end
    if (in_rt_dat_mask_d_1_46) begin
      in_rt_dat_data_d_2_46 <= in_rt_dat_data_d_1_46;
    end
    if (in_rt_dat_mask_d_1_47) begin
      in_rt_dat_data_d_2_47 <= in_rt_dat_data_d_1_47;
    end
    if (in_rt_dat_mask_d_1_48) begin
      in_rt_dat_data_d_2_48 <= in_rt_dat_data_d_1_48;
    end
    if (in_rt_dat_mask_d_1_49) begin
      in_rt_dat_data_d_2_49 <= in_rt_dat_data_d_1_49;
    end
    if (in_rt_dat_mask_d_1_50) begin
      in_rt_dat_data_d_2_50 <= in_rt_dat_data_d_1_50;
    end
    if (in_rt_dat_mask_d_1_51) begin
      in_rt_dat_data_d_2_51 <= in_rt_dat_data_d_1_51;
    end
    if (in_rt_dat_mask_d_1_52) begin
      in_rt_dat_data_d_2_52 <= in_rt_dat_data_d_1_52;
    end
    if (in_rt_dat_mask_d_1_53) begin
      in_rt_dat_data_d_2_53 <= in_rt_dat_data_d_1_53;
    end
    if (in_rt_dat_mask_d_1_54) begin
      in_rt_dat_data_d_2_54 <= in_rt_dat_data_d_1_54;
    end
    if (in_rt_dat_mask_d_1_55) begin
      in_rt_dat_data_d_2_55 <= in_rt_dat_data_d_1_55;
    end
    if (in_rt_dat_mask_d_1_56) begin
      in_rt_dat_data_d_2_56 <= in_rt_dat_data_d_1_56;
    end
    if (in_rt_dat_mask_d_1_57) begin
      in_rt_dat_data_d_2_57 <= in_rt_dat_data_d_1_57;
    end
    if (in_rt_dat_mask_d_1_58) begin
      in_rt_dat_data_d_2_58 <= in_rt_dat_data_d_1_58;
    end
    if (in_rt_dat_mask_d_1_59) begin
      in_rt_dat_data_d_2_59 <= in_rt_dat_data_d_1_59;
    end
    if (in_rt_dat_mask_d_1_60) begin
      in_rt_dat_data_d_2_60 <= in_rt_dat_data_d_1_60;
    end
    if (in_rt_dat_mask_d_1_61) begin
      in_rt_dat_data_d_2_61 <= in_rt_dat_data_d_1_61;
    end
    if (in_rt_dat_mask_d_1_62) begin
      in_rt_dat_data_d_2_62 <= in_rt_dat_data_d_1_62;
    end
    if (in_rt_dat_mask_d_1_63) begin
      in_rt_dat_data_d_2_63 <= in_rt_dat_data_d_1_63;
    end
    if (in_rt_dat_mask_d_1_64) begin
      in_rt_dat_data_d_2_64 <= in_rt_dat_data_d_1_64;
    end
    if (in_rt_dat_mask_d_1_65) begin
      in_rt_dat_data_d_2_65 <= in_rt_dat_data_d_1_65;
    end
    if (in_rt_dat_mask_d_1_66) begin
      in_rt_dat_data_d_2_66 <= in_rt_dat_data_d_1_66;
    end
    if (in_rt_dat_mask_d_1_67) begin
      in_rt_dat_data_d_2_67 <= in_rt_dat_data_d_1_67;
    end
    if (in_rt_dat_mask_d_1_68) begin
      in_rt_dat_data_d_2_68 <= in_rt_dat_data_d_1_68;
    end
    if (in_rt_dat_mask_d_1_69) begin
      in_rt_dat_data_d_2_69 <= in_rt_dat_data_d_1_69;
    end
    if (in_rt_dat_mask_d_1_70) begin
      in_rt_dat_data_d_2_70 <= in_rt_dat_data_d_1_70;
    end
    if (in_rt_dat_mask_d_1_71) begin
      in_rt_dat_data_d_2_71 <= in_rt_dat_data_d_1_71;
    end
    if (in_rt_dat_mask_d_1_72) begin
      in_rt_dat_data_d_2_72 <= in_rt_dat_data_d_1_72;
    end
    if (in_rt_dat_mask_d_1_73) begin
      in_rt_dat_data_d_2_73 <= in_rt_dat_data_d_1_73;
    end
    if (in_rt_dat_mask_d_1_74) begin
      in_rt_dat_data_d_2_74 <= in_rt_dat_data_d_1_74;
    end
    if (in_rt_dat_mask_d_1_75) begin
      in_rt_dat_data_d_2_75 <= in_rt_dat_data_d_1_75;
    end
    if (in_rt_dat_mask_d_1_76) begin
      in_rt_dat_data_d_2_76 <= in_rt_dat_data_d_1_76;
    end
    if (in_rt_dat_mask_d_1_77) begin
      in_rt_dat_data_d_2_77 <= in_rt_dat_data_d_1_77;
    end
    if (in_rt_dat_mask_d_1_78) begin
      in_rt_dat_data_d_2_78 <= in_rt_dat_data_d_1_78;
    end
    if (in_rt_dat_mask_d_1_79) begin
      in_rt_dat_data_d_2_79 <= in_rt_dat_data_d_1_79;
    end
    if (in_rt_dat_mask_d_1_80) begin
      in_rt_dat_data_d_2_80 <= in_rt_dat_data_d_1_80;
    end
    if (in_rt_dat_mask_d_1_81) begin
      in_rt_dat_data_d_2_81 <= in_rt_dat_data_d_1_81;
    end
    if (in_rt_dat_mask_d_1_82) begin
      in_rt_dat_data_d_2_82 <= in_rt_dat_data_d_1_82;
    end
    if (in_rt_dat_mask_d_1_83) begin
      in_rt_dat_data_d_2_83 <= in_rt_dat_data_d_1_83;
    end
    if (in_rt_dat_mask_d_1_84) begin
      in_rt_dat_data_d_2_84 <= in_rt_dat_data_d_1_84;
    end
    if (in_rt_dat_mask_d_1_85) begin
      in_rt_dat_data_d_2_85 <= in_rt_dat_data_d_1_85;
    end
    if (in_rt_dat_mask_d_1_86) begin
      in_rt_dat_data_d_2_86 <= in_rt_dat_data_d_1_86;
    end
    if (in_rt_dat_mask_d_1_87) begin
      in_rt_dat_data_d_2_87 <= in_rt_dat_data_d_1_87;
    end
    if (in_rt_dat_mask_d_1_88) begin
      in_rt_dat_data_d_2_88 <= in_rt_dat_data_d_1_88;
    end
    if (in_rt_dat_mask_d_1_89) begin
      in_rt_dat_data_d_2_89 <= in_rt_dat_data_d_1_89;
    end
    if (in_rt_dat_mask_d_1_90) begin
      in_rt_dat_data_d_2_90 <= in_rt_dat_data_d_1_90;
    end
    if (in_rt_dat_mask_d_1_91) begin
      in_rt_dat_data_d_2_91 <= in_rt_dat_data_d_1_91;
    end
    if (in_rt_dat_mask_d_1_92) begin
      in_rt_dat_data_d_2_92 <= in_rt_dat_data_d_1_92;
    end
    if (in_rt_dat_mask_d_1_93) begin
      in_rt_dat_data_d_2_93 <= in_rt_dat_data_d_1_93;
    end
    if (in_rt_dat_mask_d_1_94) begin
      in_rt_dat_data_d_2_94 <= in_rt_dat_data_d_1_94;
    end
    if (in_rt_dat_mask_d_1_95) begin
      in_rt_dat_data_d_2_95 <= in_rt_dat_data_d_1_95;
    end
    if (in_rt_dat_mask_d_1_96) begin
      in_rt_dat_data_d_2_96 <= in_rt_dat_data_d_1_96;
    end
    if (in_rt_dat_mask_d_1_97) begin
      in_rt_dat_data_d_2_97 <= in_rt_dat_data_d_1_97;
    end
    if (in_rt_dat_mask_d_1_98) begin
      in_rt_dat_data_d_2_98 <= in_rt_dat_data_d_1_98;
    end
    if (in_rt_dat_mask_d_1_99) begin
      in_rt_dat_data_d_2_99 <= in_rt_dat_data_d_1_99;
    end
    if (in_rt_dat_mask_d_1_100) begin
      in_rt_dat_data_d_2_100 <= in_rt_dat_data_d_1_100;
    end
    if (in_rt_dat_mask_d_1_101) begin
      in_rt_dat_data_d_2_101 <= in_rt_dat_data_d_1_101;
    end
    if (in_rt_dat_mask_d_1_102) begin
      in_rt_dat_data_d_2_102 <= in_rt_dat_data_d_1_102;
    end
    if (in_rt_dat_mask_d_1_103) begin
      in_rt_dat_data_d_2_103 <= in_rt_dat_data_d_1_103;
    end
    if (in_rt_dat_mask_d_1_104) begin
      in_rt_dat_data_d_2_104 <= in_rt_dat_data_d_1_104;
    end
    if (in_rt_dat_mask_d_1_105) begin
      in_rt_dat_data_d_2_105 <= in_rt_dat_data_d_1_105;
    end
    if (in_rt_dat_mask_d_1_106) begin
      in_rt_dat_data_d_2_106 <= in_rt_dat_data_d_1_106;
    end
    if (in_rt_dat_mask_d_1_107) begin
      in_rt_dat_data_d_2_107 <= in_rt_dat_data_d_1_107;
    end
    if (in_rt_dat_mask_d_1_108) begin
      in_rt_dat_data_d_2_108 <= in_rt_dat_data_d_1_108;
    end
    if (in_rt_dat_mask_d_1_109) begin
      in_rt_dat_data_d_2_109 <= in_rt_dat_data_d_1_109;
    end
    if (in_rt_dat_mask_d_1_110) begin
      in_rt_dat_data_d_2_110 <= in_rt_dat_data_d_1_110;
    end
    if (in_rt_dat_mask_d_1_111) begin
      in_rt_dat_data_d_2_111 <= in_rt_dat_data_d_1_111;
    end
    if (in_rt_dat_mask_d_1_112) begin
      in_rt_dat_data_d_2_112 <= in_rt_dat_data_d_1_112;
    end
    if (in_rt_dat_mask_d_1_113) begin
      in_rt_dat_data_d_2_113 <= in_rt_dat_data_d_1_113;
    end
    if (in_rt_dat_mask_d_1_114) begin
      in_rt_dat_data_d_2_114 <= in_rt_dat_data_d_1_114;
    end
    if (in_rt_dat_mask_d_1_115) begin
      in_rt_dat_data_d_2_115 <= in_rt_dat_data_d_1_115;
    end
    if (in_rt_dat_mask_d_1_116) begin
      in_rt_dat_data_d_2_116 <= in_rt_dat_data_d_1_116;
    end
    if (in_rt_dat_mask_d_1_117) begin
      in_rt_dat_data_d_2_117 <= in_rt_dat_data_d_1_117;
    end
    if (in_rt_dat_mask_d_1_118) begin
      in_rt_dat_data_d_2_118 <= in_rt_dat_data_d_1_118;
    end
    if (in_rt_dat_mask_d_1_119) begin
      in_rt_dat_data_d_2_119 <= in_rt_dat_data_d_1_119;
    end
    if (in_rt_dat_mask_d_1_120) begin
      in_rt_dat_data_d_2_120 <= in_rt_dat_data_d_1_120;
    end
    if (in_rt_dat_mask_d_1_121) begin
      in_rt_dat_data_d_2_121 <= in_rt_dat_data_d_1_121;
    end
    if (in_rt_dat_mask_d_1_122) begin
      in_rt_dat_data_d_2_122 <= in_rt_dat_data_d_1_122;
    end
    if (in_rt_dat_mask_d_1_123) begin
      in_rt_dat_data_d_2_123 <= in_rt_dat_data_d_1_123;
    end
    if (in_rt_dat_mask_d_1_124) begin
      in_rt_dat_data_d_2_124 <= in_rt_dat_data_d_1_124;
    end
    if (in_rt_dat_mask_d_1_125) begin
      in_rt_dat_data_d_2_125 <= in_rt_dat_data_d_1_125;
    end
    if (in_rt_dat_mask_d_1_126) begin
      in_rt_dat_data_d_2_126 <= in_rt_dat_data_d_1_126;
    end
    if (in_rt_dat_mask_d_1_127) begin
      in_rt_dat_data_d_2_127 <= in_rt_dat_data_d_1_127;
    end
    if (reset) begin
      in_rt_dat_mask_d_1_0 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_0 <= io_sc2mac_dat_mask_0;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_1 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_1 <= io_sc2mac_dat_mask_1;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_2 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_2 <= io_sc2mac_dat_mask_2;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_3 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_3 <= io_sc2mac_dat_mask_3;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_4 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_4 <= io_sc2mac_dat_mask_4;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_5 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_5 <= io_sc2mac_dat_mask_5;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_6 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_6 <= io_sc2mac_dat_mask_6;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_7 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_7 <= io_sc2mac_dat_mask_7;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_8 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_8 <= io_sc2mac_dat_mask_8;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_9 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_9 <= io_sc2mac_dat_mask_9;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_10 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_10 <= io_sc2mac_dat_mask_10;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_11 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_11 <= io_sc2mac_dat_mask_11;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_12 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_12 <= io_sc2mac_dat_mask_12;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_13 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_13 <= io_sc2mac_dat_mask_13;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_14 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_14 <= io_sc2mac_dat_mask_14;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_15 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_15 <= io_sc2mac_dat_mask_15;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_16 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_16 <= io_sc2mac_dat_mask_16;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_17 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_17 <= io_sc2mac_dat_mask_17;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_18 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_18 <= io_sc2mac_dat_mask_18;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_19 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_19 <= io_sc2mac_dat_mask_19;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_20 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_20 <= io_sc2mac_dat_mask_20;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_21 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_21 <= io_sc2mac_dat_mask_21;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_22 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_22 <= io_sc2mac_dat_mask_22;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_23 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_23 <= io_sc2mac_dat_mask_23;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_24 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_24 <= io_sc2mac_dat_mask_24;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_25 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_25 <= io_sc2mac_dat_mask_25;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_26 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_26 <= io_sc2mac_dat_mask_26;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_27 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_27 <= io_sc2mac_dat_mask_27;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_28 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_28 <= io_sc2mac_dat_mask_28;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_29 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_29 <= io_sc2mac_dat_mask_29;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_30 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_30 <= io_sc2mac_dat_mask_30;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_31 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_31 <= io_sc2mac_dat_mask_31;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_32 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_32 <= io_sc2mac_dat_mask_32;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_33 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_33 <= io_sc2mac_dat_mask_33;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_34 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_34 <= io_sc2mac_dat_mask_34;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_35 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_35 <= io_sc2mac_dat_mask_35;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_36 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_36 <= io_sc2mac_dat_mask_36;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_37 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_37 <= io_sc2mac_dat_mask_37;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_38 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_38 <= io_sc2mac_dat_mask_38;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_39 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_39 <= io_sc2mac_dat_mask_39;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_40 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_40 <= io_sc2mac_dat_mask_40;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_41 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_41 <= io_sc2mac_dat_mask_41;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_42 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_42 <= io_sc2mac_dat_mask_42;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_43 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_43 <= io_sc2mac_dat_mask_43;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_44 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_44 <= io_sc2mac_dat_mask_44;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_45 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_45 <= io_sc2mac_dat_mask_45;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_46 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_46 <= io_sc2mac_dat_mask_46;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_47 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_47 <= io_sc2mac_dat_mask_47;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_48 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_48 <= io_sc2mac_dat_mask_48;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_49 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_49 <= io_sc2mac_dat_mask_49;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_50 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_50 <= io_sc2mac_dat_mask_50;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_51 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_51 <= io_sc2mac_dat_mask_51;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_52 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_52 <= io_sc2mac_dat_mask_52;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_53 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_53 <= io_sc2mac_dat_mask_53;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_54 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_54 <= io_sc2mac_dat_mask_54;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_55 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_55 <= io_sc2mac_dat_mask_55;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_56 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_56 <= io_sc2mac_dat_mask_56;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_57 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_57 <= io_sc2mac_dat_mask_57;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_58 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_58 <= io_sc2mac_dat_mask_58;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_59 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_59 <= io_sc2mac_dat_mask_59;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_60 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_60 <= io_sc2mac_dat_mask_60;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_61 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_61 <= io_sc2mac_dat_mask_61;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_62 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_62 <= io_sc2mac_dat_mask_62;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_63 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_63 <= io_sc2mac_dat_mask_63;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_64 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_64 <= io_sc2mac_dat_mask_64;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_65 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_65 <= io_sc2mac_dat_mask_65;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_66 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_66 <= io_sc2mac_dat_mask_66;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_67 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_67 <= io_sc2mac_dat_mask_67;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_68 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_68 <= io_sc2mac_dat_mask_68;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_69 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_69 <= io_sc2mac_dat_mask_69;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_70 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_70 <= io_sc2mac_dat_mask_70;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_71 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_71 <= io_sc2mac_dat_mask_71;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_72 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_72 <= io_sc2mac_dat_mask_72;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_73 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_73 <= io_sc2mac_dat_mask_73;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_74 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_74 <= io_sc2mac_dat_mask_74;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_75 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_75 <= io_sc2mac_dat_mask_75;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_76 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_76 <= io_sc2mac_dat_mask_76;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_77 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_77 <= io_sc2mac_dat_mask_77;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_78 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_78 <= io_sc2mac_dat_mask_78;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_79 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_79 <= io_sc2mac_dat_mask_79;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_80 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_80 <= io_sc2mac_dat_mask_80;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_81 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_81 <= io_sc2mac_dat_mask_81;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_82 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_82 <= io_sc2mac_dat_mask_82;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_83 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_83 <= io_sc2mac_dat_mask_83;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_84 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_84 <= io_sc2mac_dat_mask_84;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_85 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_85 <= io_sc2mac_dat_mask_85;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_86 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_86 <= io_sc2mac_dat_mask_86;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_87 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_87 <= io_sc2mac_dat_mask_87;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_88 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_88 <= io_sc2mac_dat_mask_88;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_89 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_89 <= io_sc2mac_dat_mask_89;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_90 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_90 <= io_sc2mac_dat_mask_90;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_91 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_91 <= io_sc2mac_dat_mask_91;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_92 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_92 <= io_sc2mac_dat_mask_92;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_93 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_93 <= io_sc2mac_dat_mask_93;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_94 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_94 <= io_sc2mac_dat_mask_94;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_95 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_95 <= io_sc2mac_dat_mask_95;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_96 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_96 <= io_sc2mac_dat_mask_96;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_97 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_97 <= io_sc2mac_dat_mask_97;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_98 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_98 <= io_sc2mac_dat_mask_98;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_99 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_99 <= io_sc2mac_dat_mask_99;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_100 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_100 <= io_sc2mac_dat_mask_100;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_101 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_101 <= io_sc2mac_dat_mask_101;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_102 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_102 <= io_sc2mac_dat_mask_102;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_103 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_103 <= io_sc2mac_dat_mask_103;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_104 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_104 <= io_sc2mac_dat_mask_104;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_105 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_105 <= io_sc2mac_dat_mask_105;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_106 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_106 <= io_sc2mac_dat_mask_106;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_107 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_107 <= io_sc2mac_dat_mask_107;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_108 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_108 <= io_sc2mac_dat_mask_108;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_109 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_109 <= io_sc2mac_dat_mask_109;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_110 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_110 <= io_sc2mac_dat_mask_110;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_111 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_111 <= io_sc2mac_dat_mask_111;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_112 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_112 <= io_sc2mac_dat_mask_112;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_113 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_113 <= io_sc2mac_dat_mask_113;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_114 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_114 <= io_sc2mac_dat_mask_114;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_115 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_115 <= io_sc2mac_dat_mask_115;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_116 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_116 <= io_sc2mac_dat_mask_116;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_117 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_117 <= io_sc2mac_dat_mask_117;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_118 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_118 <= io_sc2mac_dat_mask_118;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_119 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_119 <= io_sc2mac_dat_mask_119;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_120 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_120 <= io_sc2mac_dat_mask_120;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_121 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_121 <= io_sc2mac_dat_mask_121;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_122 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_122 <= io_sc2mac_dat_mask_122;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_123 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_123 <= io_sc2mac_dat_mask_123;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_124 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_124 <= io_sc2mac_dat_mask_124;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_125 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_125 <= io_sc2mac_dat_mask_125;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_126 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_126 <= io_sc2mac_dat_mask_126;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_1_127 <= 1'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_mask_d_1_127 <= io_sc2mac_dat_mask_127;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_0 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_0 <= in_rt_dat_mask_d_1_0;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_1 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_1 <= in_rt_dat_mask_d_1_1;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_2 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_2 <= in_rt_dat_mask_d_1_2;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_3 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_3 <= in_rt_dat_mask_d_1_3;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_4 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_4 <= in_rt_dat_mask_d_1_4;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_5 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_5 <= in_rt_dat_mask_d_1_5;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_6 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_6 <= in_rt_dat_mask_d_1_6;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_7 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_7 <= in_rt_dat_mask_d_1_7;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_8 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_8 <= in_rt_dat_mask_d_1_8;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_9 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_9 <= in_rt_dat_mask_d_1_9;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_10 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_10 <= in_rt_dat_mask_d_1_10;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_11 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_11 <= in_rt_dat_mask_d_1_11;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_12 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_12 <= in_rt_dat_mask_d_1_12;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_13 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_13 <= in_rt_dat_mask_d_1_13;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_14 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_14 <= in_rt_dat_mask_d_1_14;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_15 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_15 <= in_rt_dat_mask_d_1_15;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_16 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_16 <= in_rt_dat_mask_d_1_16;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_17 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_17 <= in_rt_dat_mask_d_1_17;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_18 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_18 <= in_rt_dat_mask_d_1_18;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_19 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_19 <= in_rt_dat_mask_d_1_19;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_20 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_20 <= in_rt_dat_mask_d_1_20;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_21 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_21 <= in_rt_dat_mask_d_1_21;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_22 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_22 <= in_rt_dat_mask_d_1_22;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_23 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_23 <= in_rt_dat_mask_d_1_23;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_24 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_24 <= in_rt_dat_mask_d_1_24;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_25 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_25 <= in_rt_dat_mask_d_1_25;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_26 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_26 <= in_rt_dat_mask_d_1_26;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_27 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_27 <= in_rt_dat_mask_d_1_27;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_28 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_28 <= in_rt_dat_mask_d_1_28;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_29 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_29 <= in_rt_dat_mask_d_1_29;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_30 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_30 <= in_rt_dat_mask_d_1_30;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_31 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_31 <= in_rt_dat_mask_d_1_31;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_32 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_32 <= in_rt_dat_mask_d_1_32;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_33 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_33 <= in_rt_dat_mask_d_1_33;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_34 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_34 <= in_rt_dat_mask_d_1_34;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_35 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_35 <= in_rt_dat_mask_d_1_35;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_36 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_36 <= in_rt_dat_mask_d_1_36;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_37 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_37 <= in_rt_dat_mask_d_1_37;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_38 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_38 <= in_rt_dat_mask_d_1_38;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_39 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_39 <= in_rt_dat_mask_d_1_39;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_40 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_40 <= in_rt_dat_mask_d_1_40;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_41 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_41 <= in_rt_dat_mask_d_1_41;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_42 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_42 <= in_rt_dat_mask_d_1_42;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_43 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_43 <= in_rt_dat_mask_d_1_43;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_44 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_44 <= in_rt_dat_mask_d_1_44;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_45 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_45 <= in_rt_dat_mask_d_1_45;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_46 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_46 <= in_rt_dat_mask_d_1_46;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_47 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_47 <= in_rt_dat_mask_d_1_47;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_48 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_48 <= in_rt_dat_mask_d_1_48;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_49 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_49 <= in_rt_dat_mask_d_1_49;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_50 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_50 <= in_rt_dat_mask_d_1_50;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_51 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_51 <= in_rt_dat_mask_d_1_51;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_52 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_52 <= in_rt_dat_mask_d_1_52;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_53 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_53 <= in_rt_dat_mask_d_1_53;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_54 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_54 <= in_rt_dat_mask_d_1_54;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_55 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_55 <= in_rt_dat_mask_d_1_55;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_56 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_56 <= in_rt_dat_mask_d_1_56;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_57 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_57 <= in_rt_dat_mask_d_1_57;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_58 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_58 <= in_rt_dat_mask_d_1_58;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_59 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_59 <= in_rt_dat_mask_d_1_59;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_60 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_60 <= in_rt_dat_mask_d_1_60;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_61 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_61 <= in_rt_dat_mask_d_1_61;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_62 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_62 <= in_rt_dat_mask_d_1_62;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_63 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_63 <= in_rt_dat_mask_d_1_63;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_64 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_64 <= in_rt_dat_mask_d_1_64;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_65 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_65 <= in_rt_dat_mask_d_1_65;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_66 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_66 <= in_rt_dat_mask_d_1_66;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_67 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_67 <= in_rt_dat_mask_d_1_67;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_68 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_68 <= in_rt_dat_mask_d_1_68;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_69 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_69 <= in_rt_dat_mask_d_1_69;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_70 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_70 <= in_rt_dat_mask_d_1_70;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_71 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_71 <= in_rt_dat_mask_d_1_71;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_72 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_72 <= in_rt_dat_mask_d_1_72;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_73 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_73 <= in_rt_dat_mask_d_1_73;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_74 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_74 <= in_rt_dat_mask_d_1_74;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_75 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_75 <= in_rt_dat_mask_d_1_75;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_76 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_76 <= in_rt_dat_mask_d_1_76;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_77 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_77 <= in_rt_dat_mask_d_1_77;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_78 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_78 <= in_rt_dat_mask_d_1_78;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_79 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_79 <= in_rt_dat_mask_d_1_79;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_80 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_80 <= in_rt_dat_mask_d_1_80;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_81 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_81 <= in_rt_dat_mask_d_1_81;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_82 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_82 <= in_rt_dat_mask_d_1_82;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_83 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_83 <= in_rt_dat_mask_d_1_83;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_84 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_84 <= in_rt_dat_mask_d_1_84;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_85 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_85 <= in_rt_dat_mask_d_1_85;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_86 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_86 <= in_rt_dat_mask_d_1_86;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_87 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_87 <= in_rt_dat_mask_d_1_87;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_88 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_88 <= in_rt_dat_mask_d_1_88;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_89 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_89 <= in_rt_dat_mask_d_1_89;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_90 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_90 <= in_rt_dat_mask_d_1_90;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_91 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_91 <= in_rt_dat_mask_d_1_91;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_92 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_92 <= in_rt_dat_mask_d_1_92;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_93 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_93 <= in_rt_dat_mask_d_1_93;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_94 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_94 <= in_rt_dat_mask_d_1_94;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_95 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_95 <= in_rt_dat_mask_d_1_95;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_96 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_96 <= in_rt_dat_mask_d_1_96;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_97 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_97 <= in_rt_dat_mask_d_1_97;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_98 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_98 <= in_rt_dat_mask_d_1_98;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_99 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_99 <= in_rt_dat_mask_d_1_99;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_100 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_100 <= in_rt_dat_mask_d_1_100;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_101 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_101 <= in_rt_dat_mask_d_1_101;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_102 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_102 <= in_rt_dat_mask_d_1_102;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_103 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_103 <= in_rt_dat_mask_d_1_103;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_104 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_104 <= in_rt_dat_mask_d_1_104;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_105 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_105 <= in_rt_dat_mask_d_1_105;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_106 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_106 <= in_rt_dat_mask_d_1_106;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_107 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_107 <= in_rt_dat_mask_d_1_107;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_108 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_108 <= in_rt_dat_mask_d_1_108;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_109 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_109 <= in_rt_dat_mask_d_1_109;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_110 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_110 <= in_rt_dat_mask_d_1_110;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_111 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_111 <= in_rt_dat_mask_d_1_111;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_112 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_112 <= in_rt_dat_mask_d_1_112;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_113 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_113 <= in_rt_dat_mask_d_1_113;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_114 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_114 <= in_rt_dat_mask_d_1_114;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_115 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_115 <= in_rt_dat_mask_d_1_115;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_116 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_116 <= in_rt_dat_mask_d_1_116;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_117 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_117 <= in_rt_dat_mask_d_1_117;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_118 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_118 <= in_rt_dat_mask_d_1_118;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_119 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_119 <= in_rt_dat_mask_d_1_119;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_120 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_120 <= in_rt_dat_mask_d_1_120;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_121 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_121 <= in_rt_dat_mask_d_1_121;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_122 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_122 <= in_rt_dat_mask_d_1_122;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_123 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_123 <= in_rt_dat_mask_d_1_123;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_124 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_124 <= in_rt_dat_mask_d_1_124;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_125 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_125 <= in_rt_dat_mask_d_1_125;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_126 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_126 <= in_rt_dat_mask_d_1_126;
      end
    end
    if (reset) begin
      in_rt_dat_mask_d_2_127 <= 1'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_mask_d_2_127 <= in_rt_dat_mask_d_1_127;
      end
    end
    if (reset) begin
      in_rt_dat_pvld_d_1 <= 1'h0;
    end else begin
      in_rt_dat_pvld_d_1 <= io_sc2mac_dat_pvld;
    end
    if (reset) begin
      in_rt_dat_pvld_d_2 <= 1'h0;
    end else begin
      in_rt_dat_pvld_d_2 <= in_rt_dat_pvld_d_1;
    end
    if (reset) begin
      in_rt_dat_pd_d_1 <= 9'h0;
    end else begin
      if (_T_6928) begin
        in_rt_dat_pd_d_1 <= io_sc2mac_dat_pd;
      end
    end
    if (reset) begin
      in_rt_dat_pd_d_2 <= 9'h0;
    end else begin
      if (_T_6930) begin
        in_rt_dat_pd_d_2 <= in_rt_dat_pd_d_1;
      end
    end
    if (io_sc2mac_wt_mask_0) begin
      in_rt_wt_data_d_1_0 <= io_sc2mac_wt_data_0;
    end
    if (io_sc2mac_wt_mask_1) begin
      in_rt_wt_data_d_1_1 <= io_sc2mac_wt_data_1;
    end
    if (io_sc2mac_wt_mask_2) begin
      in_rt_wt_data_d_1_2 <= io_sc2mac_wt_data_2;
    end
    if (io_sc2mac_wt_mask_3) begin
      in_rt_wt_data_d_1_3 <= io_sc2mac_wt_data_3;
    end
    if (io_sc2mac_wt_mask_4) begin
      in_rt_wt_data_d_1_4 <= io_sc2mac_wt_data_4;
    end
    if (io_sc2mac_wt_mask_5) begin
      in_rt_wt_data_d_1_5 <= io_sc2mac_wt_data_5;
    end
    if (io_sc2mac_wt_mask_6) begin
      in_rt_wt_data_d_1_6 <= io_sc2mac_wt_data_6;
    end
    if (io_sc2mac_wt_mask_7) begin
      in_rt_wt_data_d_1_7 <= io_sc2mac_wt_data_7;
    end
    if (io_sc2mac_wt_mask_8) begin
      in_rt_wt_data_d_1_8 <= io_sc2mac_wt_data_8;
    end
    if (io_sc2mac_wt_mask_9) begin
      in_rt_wt_data_d_1_9 <= io_sc2mac_wt_data_9;
    end
    if (io_sc2mac_wt_mask_10) begin
      in_rt_wt_data_d_1_10 <= io_sc2mac_wt_data_10;
    end
    if (io_sc2mac_wt_mask_11) begin
      in_rt_wt_data_d_1_11 <= io_sc2mac_wt_data_11;
    end
    if (io_sc2mac_wt_mask_12) begin
      in_rt_wt_data_d_1_12 <= io_sc2mac_wt_data_12;
    end
    if (io_sc2mac_wt_mask_13) begin
      in_rt_wt_data_d_1_13 <= io_sc2mac_wt_data_13;
    end
    if (io_sc2mac_wt_mask_14) begin
      in_rt_wt_data_d_1_14 <= io_sc2mac_wt_data_14;
    end
    if (io_sc2mac_wt_mask_15) begin
      in_rt_wt_data_d_1_15 <= io_sc2mac_wt_data_15;
    end
    if (io_sc2mac_wt_mask_16) begin
      in_rt_wt_data_d_1_16 <= io_sc2mac_wt_data_16;
    end
    if (io_sc2mac_wt_mask_17) begin
      in_rt_wt_data_d_1_17 <= io_sc2mac_wt_data_17;
    end
    if (io_sc2mac_wt_mask_18) begin
      in_rt_wt_data_d_1_18 <= io_sc2mac_wt_data_18;
    end
    if (io_sc2mac_wt_mask_19) begin
      in_rt_wt_data_d_1_19 <= io_sc2mac_wt_data_19;
    end
    if (io_sc2mac_wt_mask_20) begin
      in_rt_wt_data_d_1_20 <= io_sc2mac_wt_data_20;
    end
    if (io_sc2mac_wt_mask_21) begin
      in_rt_wt_data_d_1_21 <= io_sc2mac_wt_data_21;
    end
    if (io_sc2mac_wt_mask_22) begin
      in_rt_wt_data_d_1_22 <= io_sc2mac_wt_data_22;
    end
    if (io_sc2mac_wt_mask_23) begin
      in_rt_wt_data_d_1_23 <= io_sc2mac_wt_data_23;
    end
    if (io_sc2mac_wt_mask_24) begin
      in_rt_wt_data_d_1_24 <= io_sc2mac_wt_data_24;
    end
    if (io_sc2mac_wt_mask_25) begin
      in_rt_wt_data_d_1_25 <= io_sc2mac_wt_data_25;
    end
    if (io_sc2mac_wt_mask_26) begin
      in_rt_wt_data_d_1_26 <= io_sc2mac_wt_data_26;
    end
    if (io_sc2mac_wt_mask_27) begin
      in_rt_wt_data_d_1_27 <= io_sc2mac_wt_data_27;
    end
    if (io_sc2mac_wt_mask_28) begin
      in_rt_wt_data_d_1_28 <= io_sc2mac_wt_data_28;
    end
    if (io_sc2mac_wt_mask_29) begin
      in_rt_wt_data_d_1_29 <= io_sc2mac_wt_data_29;
    end
    if (io_sc2mac_wt_mask_30) begin
      in_rt_wt_data_d_1_30 <= io_sc2mac_wt_data_30;
    end
    if (io_sc2mac_wt_mask_31) begin
      in_rt_wt_data_d_1_31 <= io_sc2mac_wt_data_31;
    end
    if (io_sc2mac_wt_mask_32) begin
      in_rt_wt_data_d_1_32 <= io_sc2mac_wt_data_32;
    end
    if (io_sc2mac_wt_mask_33) begin
      in_rt_wt_data_d_1_33 <= io_sc2mac_wt_data_33;
    end
    if (io_sc2mac_wt_mask_34) begin
      in_rt_wt_data_d_1_34 <= io_sc2mac_wt_data_34;
    end
    if (io_sc2mac_wt_mask_35) begin
      in_rt_wt_data_d_1_35 <= io_sc2mac_wt_data_35;
    end
    if (io_sc2mac_wt_mask_36) begin
      in_rt_wt_data_d_1_36 <= io_sc2mac_wt_data_36;
    end
    if (io_sc2mac_wt_mask_37) begin
      in_rt_wt_data_d_1_37 <= io_sc2mac_wt_data_37;
    end
    if (io_sc2mac_wt_mask_38) begin
      in_rt_wt_data_d_1_38 <= io_sc2mac_wt_data_38;
    end
    if (io_sc2mac_wt_mask_39) begin
      in_rt_wt_data_d_1_39 <= io_sc2mac_wt_data_39;
    end
    if (io_sc2mac_wt_mask_40) begin
      in_rt_wt_data_d_1_40 <= io_sc2mac_wt_data_40;
    end
    if (io_sc2mac_wt_mask_41) begin
      in_rt_wt_data_d_1_41 <= io_sc2mac_wt_data_41;
    end
    if (io_sc2mac_wt_mask_42) begin
      in_rt_wt_data_d_1_42 <= io_sc2mac_wt_data_42;
    end
    if (io_sc2mac_wt_mask_43) begin
      in_rt_wt_data_d_1_43 <= io_sc2mac_wt_data_43;
    end
    if (io_sc2mac_wt_mask_44) begin
      in_rt_wt_data_d_1_44 <= io_sc2mac_wt_data_44;
    end
    if (io_sc2mac_wt_mask_45) begin
      in_rt_wt_data_d_1_45 <= io_sc2mac_wt_data_45;
    end
    if (io_sc2mac_wt_mask_46) begin
      in_rt_wt_data_d_1_46 <= io_sc2mac_wt_data_46;
    end
    if (io_sc2mac_wt_mask_47) begin
      in_rt_wt_data_d_1_47 <= io_sc2mac_wt_data_47;
    end
    if (io_sc2mac_wt_mask_48) begin
      in_rt_wt_data_d_1_48 <= io_sc2mac_wt_data_48;
    end
    if (io_sc2mac_wt_mask_49) begin
      in_rt_wt_data_d_1_49 <= io_sc2mac_wt_data_49;
    end
    if (io_sc2mac_wt_mask_50) begin
      in_rt_wt_data_d_1_50 <= io_sc2mac_wt_data_50;
    end
    if (io_sc2mac_wt_mask_51) begin
      in_rt_wt_data_d_1_51 <= io_sc2mac_wt_data_51;
    end
    if (io_sc2mac_wt_mask_52) begin
      in_rt_wt_data_d_1_52 <= io_sc2mac_wt_data_52;
    end
    if (io_sc2mac_wt_mask_53) begin
      in_rt_wt_data_d_1_53 <= io_sc2mac_wt_data_53;
    end
    if (io_sc2mac_wt_mask_54) begin
      in_rt_wt_data_d_1_54 <= io_sc2mac_wt_data_54;
    end
    if (io_sc2mac_wt_mask_55) begin
      in_rt_wt_data_d_1_55 <= io_sc2mac_wt_data_55;
    end
    if (io_sc2mac_wt_mask_56) begin
      in_rt_wt_data_d_1_56 <= io_sc2mac_wt_data_56;
    end
    if (io_sc2mac_wt_mask_57) begin
      in_rt_wt_data_d_1_57 <= io_sc2mac_wt_data_57;
    end
    if (io_sc2mac_wt_mask_58) begin
      in_rt_wt_data_d_1_58 <= io_sc2mac_wt_data_58;
    end
    if (io_sc2mac_wt_mask_59) begin
      in_rt_wt_data_d_1_59 <= io_sc2mac_wt_data_59;
    end
    if (io_sc2mac_wt_mask_60) begin
      in_rt_wt_data_d_1_60 <= io_sc2mac_wt_data_60;
    end
    if (io_sc2mac_wt_mask_61) begin
      in_rt_wt_data_d_1_61 <= io_sc2mac_wt_data_61;
    end
    if (io_sc2mac_wt_mask_62) begin
      in_rt_wt_data_d_1_62 <= io_sc2mac_wt_data_62;
    end
    if (io_sc2mac_wt_mask_63) begin
      in_rt_wt_data_d_1_63 <= io_sc2mac_wt_data_63;
    end
    if (io_sc2mac_wt_mask_64) begin
      in_rt_wt_data_d_1_64 <= io_sc2mac_wt_data_64;
    end
    if (io_sc2mac_wt_mask_65) begin
      in_rt_wt_data_d_1_65 <= io_sc2mac_wt_data_65;
    end
    if (io_sc2mac_wt_mask_66) begin
      in_rt_wt_data_d_1_66 <= io_sc2mac_wt_data_66;
    end
    if (io_sc2mac_wt_mask_67) begin
      in_rt_wt_data_d_1_67 <= io_sc2mac_wt_data_67;
    end
    if (io_sc2mac_wt_mask_68) begin
      in_rt_wt_data_d_1_68 <= io_sc2mac_wt_data_68;
    end
    if (io_sc2mac_wt_mask_69) begin
      in_rt_wt_data_d_1_69 <= io_sc2mac_wt_data_69;
    end
    if (io_sc2mac_wt_mask_70) begin
      in_rt_wt_data_d_1_70 <= io_sc2mac_wt_data_70;
    end
    if (io_sc2mac_wt_mask_71) begin
      in_rt_wt_data_d_1_71 <= io_sc2mac_wt_data_71;
    end
    if (io_sc2mac_wt_mask_72) begin
      in_rt_wt_data_d_1_72 <= io_sc2mac_wt_data_72;
    end
    if (io_sc2mac_wt_mask_73) begin
      in_rt_wt_data_d_1_73 <= io_sc2mac_wt_data_73;
    end
    if (io_sc2mac_wt_mask_74) begin
      in_rt_wt_data_d_1_74 <= io_sc2mac_wt_data_74;
    end
    if (io_sc2mac_wt_mask_75) begin
      in_rt_wt_data_d_1_75 <= io_sc2mac_wt_data_75;
    end
    if (io_sc2mac_wt_mask_76) begin
      in_rt_wt_data_d_1_76 <= io_sc2mac_wt_data_76;
    end
    if (io_sc2mac_wt_mask_77) begin
      in_rt_wt_data_d_1_77 <= io_sc2mac_wt_data_77;
    end
    if (io_sc2mac_wt_mask_78) begin
      in_rt_wt_data_d_1_78 <= io_sc2mac_wt_data_78;
    end
    if (io_sc2mac_wt_mask_79) begin
      in_rt_wt_data_d_1_79 <= io_sc2mac_wt_data_79;
    end
    if (io_sc2mac_wt_mask_80) begin
      in_rt_wt_data_d_1_80 <= io_sc2mac_wt_data_80;
    end
    if (io_sc2mac_wt_mask_81) begin
      in_rt_wt_data_d_1_81 <= io_sc2mac_wt_data_81;
    end
    if (io_sc2mac_wt_mask_82) begin
      in_rt_wt_data_d_1_82 <= io_sc2mac_wt_data_82;
    end
    if (io_sc2mac_wt_mask_83) begin
      in_rt_wt_data_d_1_83 <= io_sc2mac_wt_data_83;
    end
    if (io_sc2mac_wt_mask_84) begin
      in_rt_wt_data_d_1_84 <= io_sc2mac_wt_data_84;
    end
    if (io_sc2mac_wt_mask_85) begin
      in_rt_wt_data_d_1_85 <= io_sc2mac_wt_data_85;
    end
    if (io_sc2mac_wt_mask_86) begin
      in_rt_wt_data_d_1_86 <= io_sc2mac_wt_data_86;
    end
    if (io_sc2mac_wt_mask_87) begin
      in_rt_wt_data_d_1_87 <= io_sc2mac_wt_data_87;
    end
    if (io_sc2mac_wt_mask_88) begin
      in_rt_wt_data_d_1_88 <= io_sc2mac_wt_data_88;
    end
    if (io_sc2mac_wt_mask_89) begin
      in_rt_wt_data_d_1_89 <= io_sc2mac_wt_data_89;
    end
    if (io_sc2mac_wt_mask_90) begin
      in_rt_wt_data_d_1_90 <= io_sc2mac_wt_data_90;
    end
    if (io_sc2mac_wt_mask_91) begin
      in_rt_wt_data_d_1_91 <= io_sc2mac_wt_data_91;
    end
    if (io_sc2mac_wt_mask_92) begin
      in_rt_wt_data_d_1_92 <= io_sc2mac_wt_data_92;
    end
    if (io_sc2mac_wt_mask_93) begin
      in_rt_wt_data_d_1_93 <= io_sc2mac_wt_data_93;
    end
    if (io_sc2mac_wt_mask_94) begin
      in_rt_wt_data_d_1_94 <= io_sc2mac_wt_data_94;
    end
    if (io_sc2mac_wt_mask_95) begin
      in_rt_wt_data_d_1_95 <= io_sc2mac_wt_data_95;
    end
    if (io_sc2mac_wt_mask_96) begin
      in_rt_wt_data_d_1_96 <= io_sc2mac_wt_data_96;
    end
    if (io_sc2mac_wt_mask_97) begin
      in_rt_wt_data_d_1_97 <= io_sc2mac_wt_data_97;
    end
    if (io_sc2mac_wt_mask_98) begin
      in_rt_wt_data_d_1_98 <= io_sc2mac_wt_data_98;
    end
    if (io_sc2mac_wt_mask_99) begin
      in_rt_wt_data_d_1_99 <= io_sc2mac_wt_data_99;
    end
    if (io_sc2mac_wt_mask_100) begin
      in_rt_wt_data_d_1_100 <= io_sc2mac_wt_data_100;
    end
    if (io_sc2mac_wt_mask_101) begin
      in_rt_wt_data_d_1_101 <= io_sc2mac_wt_data_101;
    end
    if (io_sc2mac_wt_mask_102) begin
      in_rt_wt_data_d_1_102 <= io_sc2mac_wt_data_102;
    end
    if (io_sc2mac_wt_mask_103) begin
      in_rt_wt_data_d_1_103 <= io_sc2mac_wt_data_103;
    end
    if (io_sc2mac_wt_mask_104) begin
      in_rt_wt_data_d_1_104 <= io_sc2mac_wt_data_104;
    end
    if (io_sc2mac_wt_mask_105) begin
      in_rt_wt_data_d_1_105 <= io_sc2mac_wt_data_105;
    end
    if (io_sc2mac_wt_mask_106) begin
      in_rt_wt_data_d_1_106 <= io_sc2mac_wt_data_106;
    end
    if (io_sc2mac_wt_mask_107) begin
      in_rt_wt_data_d_1_107 <= io_sc2mac_wt_data_107;
    end
    if (io_sc2mac_wt_mask_108) begin
      in_rt_wt_data_d_1_108 <= io_sc2mac_wt_data_108;
    end
    if (io_sc2mac_wt_mask_109) begin
      in_rt_wt_data_d_1_109 <= io_sc2mac_wt_data_109;
    end
    if (io_sc2mac_wt_mask_110) begin
      in_rt_wt_data_d_1_110 <= io_sc2mac_wt_data_110;
    end
    if (io_sc2mac_wt_mask_111) begin
      in_rt_wt_data_d_1_111 <= io_sc2mac_wt_data_111;
    end
    if (io_sc2mac_wt_mask_112) begin
      in_rt_wt_data_d_1_112 <= io_sc2mac_wt_data_112;
    end
    if (io_sc2mac_wt_mask_113) begin
      in_rt_wt_data_d_1_113 <= io_sc2mac_wt_data_113;
    end
    if (io_sc2mac_wt_mask_114) begin
      in_rt_wt_data_d_1_114 <= io_sc2mac_wt_data_114;
    end
    if (io_sc2mac_wt_mask_115) begin
      in_rt_wt_data_d_1_115 <= io_sc2mac_wt_data_115;
    end
    if (io_sc2mac_wt_mask_116) begin
      in_rt_wt_data_d_1_116 <= io_sc2mac_wt_data_116;
    end
    if (io_sc2mac_wt_mask_117) begin
      in_rt_wt_data_d_1_117 <= io_sc2mac_wt_data_117;
    end
    if (io_sc2mac_wt_mask_118) begin
      in_rt_wt_data_d_1_118 <= io_sc2mac_wt_data_118;
    end
    if (io_sc2mac_wt_mask_119) begin
      in_rt_wt_data_d_1_119 <= io_sc2mac_wt_data_119;
    end
    if (io_sc2mac_wt_mask_120) begin
      in_rt_wt_data_d_1_120 <= io_sc2mac_wt_data_120;
    end
    if (io_sc2mac_wt_mask_121) begin
      in_rt_wt_data_d_1_121 <= io_sc2mac_wt_data_121;
    end
    if (io_sc2mac_wt_mask_122) begin
      in_rt_wt_data_d_1_122 <= io_sc2mac_wt_data_122;
    end
    if (io_sc2mac_wt_mask_123) begin
      in_rt_wt_data_d_1_123 <= io_sc2mac_wt_data_123;
    end
    if (io_sc2mac_wt_mask_124) begin
      in_rt_wt_data_d_1_124 <= io_sc2mac_wt_data_124;
    end
    if (io_sc2mac_wt_mask_125) begin
      in_rt_wt_data_d_1_125 <= io_sc2mac_wt_data_125;
    end
    if (io_sc2mac_wt_mask_126) begin
      in_rt_wt_data_d_1_126 <= io_sc2mac_wt_data_126;
    end
    if (io_sc2mac_wt_mask_127) begin
      in_rt_wt_data_d_1_127 <= io_sc2mac_wt_data_127;
    end
    if (in_rt_wt_mask_d_1_0) begin
      in_rt_wt_data_d_2_0 <= in_rt_wt_data_d_1_0;
    end
    if (in_rt_wt_mask_d_1_1) begin
      in_rt_wt_data_d_2_1 <= in_rt_wt_data_d_1_1;
    end
    if (in_rt_wt_mask_d_1_2) begin
      in_rt_wt_data_d_2_2 <= in_rt_wt_data_d_1_2;
    end
    if (in_rt_wt_mask_d_1_3) begin
      in_rt_wt_data_d_2_3 <= in_rt_wt_data_d_1_3;
    end
    if (in_rt_wt_mask_d_1_4) begin
      in_rt_wt_data_d_2_4 <= in_rt_wt_data_d_1_4;
    end
    if (in_rt_wt_mask_d_1_5) begin
      in_rt_wt_data_d_2_5 <= in_rt_wt_data_d_1_5;
    end
    if (in_rt_wt_mask_d_1_6) begin
      in_rt_wt_data_d_2_6 <= in_rt_wt_data_d_1_6;
    end
    if (in_rt_wt_mask_d_1_7) begin
      in_rt_wt_data_d_2_7 <= in_rt_wt_data_d_1_7;
    end
    if (in_rt_wt_mask_d_1_8) begin
      in_rt_wt_data_d_2_8 <= in_rt_wt_data_d_1_8;
    end
    if (in_rt_wt_mask_d_1_9) begin
      in_rt_wt_data_d_2_9 <= in_rt_wt_data_d_1_9;
    end
    if (in_rt_wt_mask_d_1_10) begin
      in_rt_wt_data_d_2_10 <= in_rt_wt_data_d_1_10;
    end
    if (in_rt_wt_mask_d_1_11) begin
      in_rt_wt_data_d_2_11 <= in_rt_wt_data_d_1_11;
    end
    if (in_rt_wt_mask_d_1_12) begin
      in_rt_wt_data_d_2_12 <= in_rt_wt_data_d_1_12;
    end
    if (in_rt_wt_mask_d_1_13) begin
      in_rt_wt_data_d_2_13 <= in_rt_wt_data_d_1_13;
    end
    if (in_rt_wt_mask_d_1_14) begin
      in_rt_wt_data_d_2_14 <= in_rt_wt_data_d_1_14;
    end
    if (in_rt_wt_mask_d_1_15) begin
      in_rt_wt_data_d_2_15 <= in_rt_wt_data_d_1_15;
    end
    if (in_rt_wt_mask_d_1_16) begin
      in_rt_wt_data_d_2_16 <= in_rt_wt_data_d_1_16;
    end
    if (in_rt_wt_mask_d_1_17) begin
      in_rt_wt_data_d_2_17 <= in_rt_wt_data_d_1_17;
    end
    if (in_rt_wt_mask_d_1_18) begin
      in_rt_wt_data_d_2_18 <= in_rt_wt_data_d_1_18;
    end
    if (in_rt_wt_mask_d_1_19) begin
      in_rt_wt_data_d_2_19 <= in_rt_wt_data_d_1_19;
    end
    if (in_rt_wt_mask_d_1_20) begin
      in_rt_wt_data_d_2_20 <= in_rt_wt_data_d_1_20;
    end
    if (in_rt_wt_mask_d_1_21) begin
      in_rt_wt_data_d_2_21 <= in_rt_wt_data_d_1_21;
    end
    if (in_rt_wt_mask_d_1_22) begin
      in_rt_wt_data_d_2_22 <= in_rt_wt_data_d_1_22;
    end
    if (in_rt_wt_mask_d_1_23) begin
      in_rt_wt_data_d_2_23 <= in_rt_wt_data_d_1_23;
    end
    if (in_rt_wt_mask_d_1_24) begin
      in_rt_wt_data_d_2_24 <= in_rt_wt_data_d_1_24;
    end
    if (in_rt_wt_mask_d_1_25) begin
      in_rt_wt_data_d_2_25 <= in_rt_wt_data_d_1_25;
    end
    if (in_rt_wt_mask_d_1_26) begin
      in_rt_wt_data_d_2_26 <= in_rt_wt_data_d_1_26;
    end
    if (in_rt_wt_mask_d_1_27) begin
      in_rt_wt_data_d_2_27 <= in_rt_wt_data_d_1_27;
    end
    if (in_rt_wt_mask_d_1_28) begin
      in_rt_wt_data_d_2_28 <= in_rt_wt_data_d_1_28;
    end
    if (in_rt_wt_mask_d_1_29) begin
      in_rt_wt_data_d_2_29 <= in_rt_wt_data_d_1_29;
    end
    if (in_rt_wt_mask_d_1_30) begin
      in_rt_wt_data_d_2_30 <= in_rt_wt_data_d_1_30;
    end
    if (in_rt_wt_mask_d_1_31) begin
      in_rt_wt_data_d_2_31 <= in_rt_wt_data_d_1_31;
    end
    if (in_rt_wt_mask_d_1_32) begin
      in_rt_wt_data_d_2_32 <= in_rt_wt_data_d_1_32;
    end
    if (in_rt_wt_mask_d_1_33) begin
      in_rt_wt_data_d_2_33 <= in_rt_wt_data_d_1_33;
    end
    if (in_rt_wt_mask_d_1_34) begin
      in_rt_wt_data_d_2_34 <= in_rt_wt_data_d_1_34;
    end
    if (in_rt_wt_mask_d_1_35) begin
      in_rt_wt_data_d_2_35 <= in_rt_wt_data_d_1_35;
    end
    if (in_rt_wt_mask_d_1_36) begin
      in_rt_wt_data_d_2_36 <= in_rt_wt_data_d_1_36;
    end
    if (in_rt_wt_mask_d_1_37) begin
      in_rt_wt_data_d_2_37 <= in_rt_wt_data_d_1_37;
    end
    if (in_rt_wt_mask_d_1_38) begin
      in_rt_wt_data_d_2_38 <= in_rt_wt_data_d_1_38;
    end
    if (in_rt_wt_mask_d_1_39) begin
      in_rt_wt_data_d_2_39 <= in_rt_wt_data_d_1_39;
    end
    if (in_rt_wt_mask_d_1_40) begin
      in_rt_wt_data_d_2_40 <= in_rt_wt_data_d_1_40;
    end
    if (in_rt_wt_mask_d_1_41) begin
      in_rt_wt_data_d_2_41 <= in_rt_wt_data_d_1_41;
    end
    if (in_rt_wt_mask_d_1_42) begin
      in_rt_wt_data_d_2_42 <= in_rt_wt_data_d_1_42;
    end
    if (in_rt_wt_mask_d_1_43) begin
      in_rt_wt_data_d_2_43 <= in_rt_wt_data_d_1_43;
    end
    if (in_rt_wt_mask_d_1_44) begin
      in_rt_wt_data_d_2_44 <= in_rt_wt_data_d_1_44;
    end
    if (in_rt_wt_mask_d_1_45) begin
      in_rt_wt_data_d_2_45 <= in_rt_wt_data_d_1_45;
    end
    if (in_rt_wt_mask_d_1_46) begin
      in_rt_wt_data_d_2_46 <= in_rt_wt_data_d_1_46;
    end
    if (in_rt_wt_mask_d_1_47) begin
      in_rt_wt_data_d_2_47 <= in_rt_wt_data_d_1_47;
    end
    if (in_rt_wt_mask_d_1_48) begin
      in_rt_wt_data_d_2_48 <= in_rt_wt_data_d_1_48;
    end
    if (in_rt_wt_mask_d_1_49) begin
      in_rt_wt_data_d_2_49 <= in_rt_wt_data_d_1_49;
    end
    if (in_rt_wt_mask_d_1_50) begin
      in_rt_wt_data_d_2_50 <= in_rt_wt_data_d_1_50;
    end
    if (in_rt_wt_mask_d_1_51) begin
      in_rt_wt_data_d_2_51 <= in_rt_wt_data_d_1_51;
    end
    if (in_rt_wt_mask_d_1_52) begin
      in_rt_wt_data_d_2_52 <= in_rt_wt_data_d_1_52;
    end
    if (in_rt_wt_mask_d_1_53) begin
      in_rt_wt_data_d_2_53 <= in_rt_wt_data_d_1_53;
    end
    if (in_rt_wt_mask_d_1_54) begin
      in_rt_wt_data_d_2_54 <= in_rt_wt_data_d_1_54;
    end
    if (in_rt_wt_mask_d_1_55) begin
      in_rt_wt_data_d_2_55 <= in_rt_wt_data_d_1_55;
    end
    if (in_rt_wt_mask_d_1_56) begin
      in_rt_wt_data_d_2_56 <= in_rt_wt_data_d_1_56;
    end
    if (in_rt_wt_mask_d_1_57) begin
      in_rt_wt_data_d_2_57 <= in_rt_wt_data_d_1_57;
    end
    if (in_rt_wt_mask_d_1_58) begin
      in_rt_wt_data_d_2_58 <= in_rt_wt_data_d_1_58;
    end
    if (in_rt_wt_mask_d_1_59) begin
      in_rt_wt_data_d_2_59 <= in_rt_wt_data_d_1_59;
    end
    if (in_rt_wt_mask_d_1_60) begin
      in_rt_wt_data_d_2_60 <= in_rt_wt_data_d_1_60;
    end
    if (in_rt_wt_mask_d_1_61) begin
      in_rt_wt_data_d_2_61 <= in_rt_wt_data_d_1_61;
    end
    if (in_rt_wt_mask_d_1_62) begin
      in_rt_wt_data_d_2_62 <= in_rt_wt_data_d_1_62;
    end
    if (in_rt_wt_mask_d_1_63) begin
      in_rt_wt_data_d_2_63 <= in_rt_wt_data_d_1_63;
    end
    if (in_rt_wt_mask_d_1_64) begin
      in_rt_wt_data_d_2_64 <= in_rt_wt_data_d_1_64;
    end
    if (in_rt_wt_mask_d_1_65) begin
      in_rt_wt_data_d_2_65 <= in_rt_wt_data_d_1_65;
    end
    if (in_rt_wt_mask_d_1_66) begin
      in_rt_wt_data_d_2_66 <= in_rt_wt_data_d_1_66;
    end
    if (in_rt_wt_mask_d_1_67) begin
      in_rt_wt_data_d_2_67 <= in_rt_wt_data_d_1_67;
    end
    if (in_rt_wt_mask_d_1_68) begin
      in_rt_wt_data_d_2_68 <= in_rt_wt_data_d_1_68;
    end
    if (in_rt_wt_mask_d_1_69) begin
      in_rt_wt_data_d_2_69 <= in_rt_wt_data_d_1_69;
    end
    if (in_rt_wt_mask_d_1_70) begin
      in_rt_wt_data_d_2_70 <= in_rt_wt_data_d_1_70;
    end
    if (in_rt_wt_mask_d_1_71) begin
      in_rt_wt_data_d_2_71 <= in_rt_wt_data_d_1_71;
    end
    if (in_rt_wt_mask_d_1_72) begin
      in_rt_wt_data_d_2_72 <= in_rt_wt_data_d_1_72;
    end
    if (in_rt_wt_mask_d_1_73) begin
      in_rt_wt_data_d_2_73 <= in_rt_wt_data_d_1_73;
    end
    if (in_rt_wt_mask_d_1_74) begin
      in_rt_wt_data_d_2_74 <= in_rt_wt_data_d_1_74;
    end
    if (in_rt_wt_mask_d_1_75) begin
      in_rt_wt_data_d_2_75 <= in_rt_wt_data_d_1_75;
    end
    if (in_rt_wt_mask_d_1_76) begin
      in_rt_wt_data_d_2_76 <= in_rt_wt_data_d_1_76;
    end
    if (in_rt_wt_mask_d_1_77) begin
      in_rt_wt_data_d_2_77 <= in_rt_wt_data_d_1_77;
    end
    if (in_rt_wt_mask_d_1_78) begin
      in_rt_wt_data_d_2_78 <= in_rt_wt_data_d_1_78;
    end
    if (in_rt_wt_mask_d_1_79) begin
      in_rt_wt_data_d_2_79 <= in_rt_wt_data_d_1_79;
    end
    if (in_rt_wt_mask_d_1_80) begin
      in_rt_wt_data_d_2_80 <= in_rt_wt_data_d_1_80;
    end
    if (in_rt_wt_mask_d_1_81) begin
      in_rt_wt_data_d_2_81 <= in_rt_wt_data_d_1_81;
    end
    if (in_rt_wt_mask_d_1_82) begin
      in_rt_wt_data_d_2_82 <= in_rt_wt_data_d_1_82;
    end
    if (in_rt_wt_mask_d_1_83) begin
      in_rt_wt_data_d_2_83 <= in_rt_wt_data_d_1_83;
    end
    if (in_rt_wt_mask_d_1_84) begin
      in_rt_wt_data_d_2_84 <= in_rt_wt_data_d_1_84;
    end
    if (in_rt_wt_mask_d_1_85) begin
      in_rt_wt_data_d_2_85 <= in_rt_wt_data_d_1_85;
    end
    if (in_rt_wt_mask_d_1_86) begin
      in_rt_wt_data_d_2_86 <= in_rt_wt_data_d_1_86;
    end
    if (in_rt_wt_mask_d_1_87) begin
      in_rt_wt_data_d_2_87 <= in_rt_wt_data_d_1_87;
    end
    if (in_rt_wt_mask_d_1_88) begin
      in_rt_wt_data_d_2_88 <= in_rt_wt_data_d_1_88;
    end
    if (in_rt_wt_mask_d_1_89) begin
      in_rt_wt_data_d_2_89 <= in_rt_wt_data_d_1_89;
    end
    if (in_rt_wt_mask_d_1_90) begin
      in_rt_wt_data_d_2_90 <= in_rt_wt_data_d_1_90;
    end
    if (in_rt_wt_mask_d_1_91) begin
      in_rt_wt_data_d_2_91 <= in_rt_wt_data_d_1_91;
    end
    if (in_rt_wt_mask_d_1_92) begin
      in_rt_wt_data_d_2_92 <= in_rt_wt_data_d_1_92;
    end
    if (in_rt_wt_mask_d_1_93) begin
      in_rt_wt_data_d_2_93 <= in_rt_wt_data_d_1_93;
    end
    if (in_rt_wt_mask_d_1_94) begin
      in_rt_wt_data_d_2_94 <= in_rt_wt_data_d_1_94;
    end
    if (in_rt_wt_mask_d_1_95) begin
      in_rt_wt_data_d_2_95 <= in_rt_wt_data_d_1_95;
    end
    if (in_rt_wt_mask_d_1_96) begin
      in_rt_wt_data_d_2_96 <= in_rt_wt_data_d_1_96;
    end
    if (in_rt_wt_mask_d_1_97) begin
      in_rt_wt_data_d_2_97 <= in_rt_wt_data_d_1_97;
    end
    if (in_rt_wt_mask_d_1_98) begin
      in_rt_wt_data_d_2_98 <= in_rt_wt_data_d_1_98;
    end
    if (in_rt_wt_mask_d_1_99) begin
      in_rt_wt_data_d_2_99 <= in_rt_wt_data_d_1_99;
    end
    if (in_rt_wt_mask_d_1_100) begin
      in_rt_wt_data_d_2_100 <= in_rt_wt_data_d_1_100;
    end
    if (in_rt_wt_mask_d_1_101) begin
      in_rt_wt_data_d_2_101 <= in_rt_wt_data_d_1_101;
    end
    if (in_rt_wt_mask_d_1_102) begin
      in_rt_wt_data_d_2_102 <= in_rt_wt_data_d_1_102;
    end
    if (in_rt_wt_mask_d_1_103) begin
      in_rt_wt_data_d_2_103 <= in_rt_wt_data_d_1_103;
    end
    if (in_rt_wt_mask_d_1_104) begin
      in_rt_wt_data_d_2_104 <= in_rt_wt_data_d_1_104;
    end
    if (in_rt_wt_mask_d_1_105) begin
      in_rt_wt_data_d_2_105 <= in_rt_wt_data_d_1_105;
    end
    if (in_rt_wt_mask_d_1_106) begin
      in_rt_wt_data_d_2_106 <= in_rt_wt_data_d_1_106;
    end
    if (in_rt_wt_mask_d_1_107) begin
      in_rt_wt_data_d_2_107 <= in_rt_wt_data_d_1_107;
    end
    if (in_rt_wt_mask_d_1_108) begin
      in_rt_wt_data_d_2_108 <= in_rt_wt_data_d_1_108;
    end
    if (in_rt_wt_mask_d_1_109) begin
      in_rt_wt_data_d_2_109 <= in_rt_wt_data_d_1_109;
    end
    if (in_rt_wt_mask_d_1_110) begin
      in_rt_wt_data_d_2_110 <= in_rt_wt_data_d_1_110;
    end
    if (in_rt_wt_mask_d_1_111) begin
      in_rt_wt_data_d_2_111 <= in_rt_wt_data_d_1_111;
    end
    if (in_rt_wt_mask_d_1_112) begin
      in_rt_wt_data_d_2_112 <= in_rt_wt_data_d_1_112;
    end
    if (in_rt_wt_mask_d_1_113) begin
      in_rt_wt_data_d_2_113 <= in_rt_wt_data_d_1_113;
    end
    if (in_rt_wt_mask_d_1_114) begin
      in_rt_wt_data_d_2_114 <= in_rt_wt_data_d_1_114;
    end
    if (in_rt_wt_mask_d_1_115) begin
      in_rt_wt_data_d_2_115 <= in_rt_wt_data_d_1_115;
    end
    if (in_rt_wt_mask_d_1_116) begin
      in_rt_wt_data_d_2_116 <= in_rt_wt_data_d_1_116;
    end
    if (in_rt_wt_mask_d_1_117) begin
      in_rt_wt_data_d_2_117 <= in_rt_wt_data_d_1_117;
    end
    if (in_rt_wt_mask_d_1_118) begin
      in_rt_wt_data_d_2_118 <= in_rt_wt_data_d_1_118;
    end
    if (in_rt_wt_mask_d_1_119) begin
      in_rt_wt_data_d_2_119 <= in_rt_wt_data_d_1_119;
    end
    if (in_rt_wt_mask_d_1_120) begin
      in_rt_wt_data_d_2_120 <= in_rt_wt_data_d_1_120;
    end
    if (in_rt_wt_mask_d_1_121) begin
      in_rt_wt_data_d_2_121 <= in_rt_wt_data_d_1_121;
    end
    if (in_rt_wt_mask_d_1_122) begin
      in_rt_wt_data_d_2_122 <= in_rt_wt_data_d_1_122;
    end
    if (in_rt_wt_mask_d_1_123) begin
      in_rt_wt_data_d_2_123 <= in_rt_wt_data_d_1_123;
    end
    if (in_rt_wt_mask_d_1_124) begin
      in_rt_wt_data_d_2_124 <= in_rt_wt_data_d_1_124;
    end
    if (in_rt_wt_mask_d_1_125) begin
      in_rt_wt_data_d_2_125 <= in_rt_wt_data_d_1_125;
    end
    if (in_rt_wt_mask_d_1_126) begin
      in_rt_wt_data_d_2_126 <= in_rt_wt_data_d_1_126;
    end
    if (in_rt_wt_mask_d_1_127) begin
      in_rt_wt_data_d_2_127 <= in_rt_wt_data_d_1_127;
    end
    if (reset) begin
      in_rt_wt_mask_d_1_0 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_0 <= io_sc2mac_wt_mask_0;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_1 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_1 <= io_sc2mac_wt_mask_1;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_2 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_2 <= io_sc2mac_wt_mask_2;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_3 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_3 <= io_sc2mac_wt_mask_3;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_4 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_4 <= io_sc2mac_wt_mask_4;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_5 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_5 <= io_sc2mac_wt_mask_5;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_6 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_6 <= io_sc2mac_wt_mask_6;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_7 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_7 <= io_sc2mac_wt_mask_7;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_8 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_8 <= io_sc2mac_wt_mask_8;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_9 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_9 <= io_sc2mac_wt_mask_9;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_10 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_10 <= io_sc2mac_wt_mask_10;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_11 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_11 <= io_sc2mac_wt_mask_11;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_12 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_12 <= io_sc2mac_wt_mask_12;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_13 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_13 <= io_sc2mac_wt_mask_13;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_14 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_14 <= io_sc2mac_wt_mask_14;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_15 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_15 <= io_sc2mac_wt_mask_15;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_16 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_16 <= io_sc2mac_wt_mask_16;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_17 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_17 <= io_sc2mac_wt_mask_17;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_18 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_18 <= io_sc2mac_wt_mask_18;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_19 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_19 <= io_sc2mac_wt_mask_19;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_20 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_20 <= io_sc2mac_wt_mask_20;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_21 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_21 <= io_sc2mac_wt_mask_21;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_22 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_22 <= io_sc2mac_wt_mask_22;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_23 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_23 <= io_sc2mac_wt_mask_23;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_24 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_24 <= io_sc2mac_wt_mask_24;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_25 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_25 <= io_sc2mac_wt_mask_25;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_26 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_26 <= io_sc2mac_wt_mask_26;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_27 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_27 <= io_sc2mac_wt_mask_27;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_28 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_28 <= io_sc2mac_wt_mask_28;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_29 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_29 <= io_sc2mac_wt_mask_29;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_30 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_30 <= io_sc2mac_wt_mask_30;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_31 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_31 <= io_sc2mac_wt_mask_31;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_32 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_32 <= io_sc2mac_wt_mask_32;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_33 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_33 <= io_sc2mac_wt_mask_33;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_34 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_34 <= io_sc2mac_wt_mask_34;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_35 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_35 <= io_sc2mac_wt_mask_35;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_36 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_36 <= io_sc2mac_wt_mask_36;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_37 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_37 <= io_sc2mac_wt_mask_37;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_38 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_38 <= io_sc2mac_wt_mask_38;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_39 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_39 <= io_sc2mac_wt_mask_39;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_40 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_40 <= io_sc2mac_wt_mask_40;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_41 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_41 <= io_sc2mac_wt_mask_41;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_42 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_42 <= io_sc2mac_wt_mask_42;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_43 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_43 <= io_sc2mac_wt_mask_43;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_44 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_44 <= io_sc2mac_wt_mask_44;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_45 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_45 <= io_sc2mac_wt_mask_45;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_46 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_46 <= io_sc2mac_wt_mask_46;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_47 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_47 <= io_sc2mac_wt_mask_47;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_48 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_48 <= io_sc2mac_wt_mask_48;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_49 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_49 <= io_sc2mac_wt_mask_49;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_50 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_50 <= io_sc2mac_wt_mask_50;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_51 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_51 <= io_sc2mac_wt_mask_51;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_52 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_52 <= io_sc2mac_wt_mask_52;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_53 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_53 <= io_sc2mac_wt_mask_53;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_54 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_54 <= io_sc2mac_wt_mask_54;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_55 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_55 <= io_sc2mac_wt_mask_55;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_56 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_56 <= io_sc2mac_wt_mask_56;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_57 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_57 <= io_sc2mac_wt_mask_57;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_58 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_58 <= io_sc2mac_wt_mask_58;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_59 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_59 <= io_sc2mac_wt_mask_59;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_60 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_60 <= io_sc2mac_wt_mask_60;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_61 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_61 <= io_sc2mac_wt_mask_61;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_62 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_62 <= io_sc2mac_wt_mask_62;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_63 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_63 <= io_sc2mac_wt_mask_63;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_64 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_64 <= io_sc2mac_wt_mask_64;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_65 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_65 <= io_sc2mac_wt_mask_65;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_66 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_66 <= io_sc2mac_wt_mask_66;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_67 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_67 <= io_sc2mac_wt_mask_67;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_68 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_68 <= io_sc2mac_wt_mask_68;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_69 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_69 <= io_sc2mac_wt_mask_69;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_70 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_70 <= io_sc2mac_wt_mask_70;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_71 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_71 <= io_sc2mac_wt_mask_71;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_72 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_72 <= io_sc2mac_wt_mask_72;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_73 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_73 <= io_sc2mac_wt_mask_73;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_74 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_74 <= io_sc2mac_wt_mask_74;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_75 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_75 <= io_sc2mac_wt_mask_75;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_76 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_76 <= io_sc2mac_wt_mask_76;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_77 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_77 <= io_sc2mac_wt_mask_77;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_78 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_78 <= io_sc2mac_wt_mask_78;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_79 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_79 <= io_sc2mac_wt_mask_79;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_80 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_80 <= io_sc2mac_wt_mask_80;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_81 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_81 <= io_sc2mac_wt_mask_81;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_82 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_82 <= io_sc2mac_wt_mask_82;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_83 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_83 <= io_sc2mac_wt_mask_83;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_84 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_84 <= io_sc2mac_wt_mask_84;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_85 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_85 <= io_sc2mac_wt_mask_85;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_86 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_86 <= io_sc2mac_wt_mask_86;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_87 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_87 <= io_sc2mac_wt_mask_87;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_88 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_88 <= io_sc2mac_wt_mask_88;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_89 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_89 <= io_sc2mac_wt_mask_89;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_90 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_90 <= io_sc2mac_wt_mask_90;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_91 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_91 <= io_sc2mac_wt_mask_91;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_92 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_92 <= io_sc2mac_wt_mask_92;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_93 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_93 <= io_sc2mac_wt_mask_93;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_94 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_94 <= io_sc2mac_wt_mask_94;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_95 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_95 <= io_sc2mac_wt_mask_95;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_96 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_96 <= io_sc2mac_wt_mask_96;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_97 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_97 <= io_sc2mac_wt_mask_97;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_98 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_98 <= io_sc2mac_wt_mask_98;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_99 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_99 <= io_sc2mac_wt_mask_99;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_100 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_100 <= io_sc2mac_wt_mask_100;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_101 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_101 <= io_sc2mac_wt_mask_101;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_102 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_102 <= io_sc2mac_wt_mask_102;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_103 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_103 <= io_sc2mac_wt_mask_103;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_104 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_104 <= io_sc2mac_wt_mask_104;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_105 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_105 <= io_sc2mac_wt_mask_105;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_106 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_106 <= io_sc2mac_wt_mask_106;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_107 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_107 <= io_sc2mac_wt_mask_107;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_108 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_108 <= io_sc2mac_wt_mask_108;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_109 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_109 <= io_sc2mac_wt_mask_109;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_110 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_110 <= io_sc2mac_wt_mask_110;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_111 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_111 <= io_sc2mac_wt_mask_111;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_112 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_112 <= io_sc2mac_wt_mask_112;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_113 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_113 <= io_sc2mac_wt_mask_113;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_114 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_114 <= io_sc2mac_wt_mask_114;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_115 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_115 <= io_sc2mac_wt_mask_115;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_116 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_116 <= io_sc2mac_wt_mask_116;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_117 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_117 <= io_sc2mac_wt_mask_117;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_118 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_118 <= io_sc2mac_wt_mask_118;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_119 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_119 <= io_sc2mac_wt_mask_119;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_120 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_120 <= io_sc2mac_wt_mask_120;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_121 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_121 <= io_sc2mac_wt_mask_121;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_122 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_122 <= io_sc2mac_wt_mask_122;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_123 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_123 <= io_sc2mac_wt_mask_123;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_124 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_124 <= io_sc2mac_wt_mask_124;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_125 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_125 <= io_sc2mac_wt_mask_125;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_126 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_126 <= io_sc2mac_wt_mask_126;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_1_127 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_mask_d_1_127 <= io_sc2mac_wt_mask_127;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_0 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_0 <= in_rt_wt_mask_d_1_0;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_1 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_1 <= in_rt_wt_mask_d_1_1;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_2 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_2 <= in_rt_wt_mask_d_1_2;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_3 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_3 <= in_rt_wt_mask_d_1_3;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_4 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_4 <= in_rt_wt_mask_d_1_4;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_5 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_5 <= in_rt_wt_mask_d_1_5;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_6 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_6 <= in_rt_wt_mask_d_1_6;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_7 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_7 <= in_rt_wt_mask_d_1_7;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_8 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_8 <= in_rt_wt_mask_d_1_8;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_9 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_9 <= in_rt_wt_mask_d_1_9;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_10 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_10 <= in_rt_wt_mask_d_1_10;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_11 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_11 <= in_rt_wt_mask_d_1_11;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_12 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_12 <= in_rt_wt_mask_d_1_12;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_13 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_13 <= in_rt_wt_mask_d_1_13;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_14 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_14 <= in_rt_wt_mask_d_1_14;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_15 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_15 <= in_rt_wt_mask_d_1_15;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_16 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_16 <= in_rt_wt_mask_d_1_16;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_17 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_17 <= in_rt_wt_mask_d_1_17;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_18 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_18 <= in_rt_wt_mask_d_1_18;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_19 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_19 <= in_rt_wt_mask_d_1_19;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_20 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_20 <= in_rt_wt_mask_d_1_20;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_21 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_21 <= in_rt_wt_mask_d_1_21;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_22 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_22 <= in_rt_wt_mask_d_1_22;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_23 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_23 <= in_rt_wt_mask_d_1_23;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_24 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_24 <= in_rt_wt_mask_d_1_24;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_25 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_25 <= in_rt_wt_mask_d_1_25;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_26 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_26 <= in_rt_wt_mask_d_1_26;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_27 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_27 <= in_rt_wt_mask_d_1_27;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_28 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_28 <= in_rt_wt_mask_d_1_28;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_29 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_29 <= in_rt_wt_mask_d_1_29;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_30 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_30 <= in_rt_wt_mask_d_1_30;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_31 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_31 <= in_rt_wt_mask_d_1_31;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_32 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_32 <= in_rt_wt_mask_d_1_32;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_33 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_33 <= in_rt_wt_mask_d_1_33;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_34 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_34 <= in_rt_wt_mask_d_1_34;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_35 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_35 <= in_rt_wt_mask_d_1_35;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_36 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_36 <= in_rt_wt_mask_d_1_36;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_37 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_37 <= in_rt_wt_mask_d_1_37;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_38 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_38 <= in_rt_wt_mask_d_1_38;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_39 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_39 <= in_rt_wt_mask_d_1_39;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_40 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_40 <= in_rt_wt_mask_d_1_40;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_41 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_41 <= in_rt_wt_mask_d_1_41;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_42 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_42 <= in_rt_wt_mask_d_1_42;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_43 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_43 <= in_rt_wt_mask_d_1_43;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_44 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_44 <= in_rt_wt_mask_d_1_44;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_45 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_45 <= in_rt_wt_mask_d_1_45;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_46 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_46 <= in_rt_wt_mask_d_1_46;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_47 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_47 <= in_rt_wt_mask_d_1_47;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_48 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_48 <= in_rt_wt_mask_d_1_48;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_49 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_49 <= in_rt_wt_mask_d_1_49;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_50 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_50 <= in_rt_wt_mask_d_1_50;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_51 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_51 <= in_rt_wt_mask_d_1_51;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_52 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_52 <= in_rt_wt_mask_d_1_52;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_53 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_53 <= in_rt_wt_mask_d_1_53;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_54 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_54 <= in_rt_wt_mask_d_1_54;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_55 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_55 <= in_rt_wt_mask_d_1_55;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_56 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_56 <= in_rt_wt_mask_d_1_56;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_57 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_57 <= in_rt_wt_mask_d_1_57;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_58 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_58 <= in_rt_wt_mask_d_1_58;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_59 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_59 <= in_rt_wt_mask_d_1_59;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_60 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_60 <= in_rt_wt_mask_d_1_60;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_61 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_61 <= in_rt_wt_mask_d_1_61;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_62 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_62 <= in_rt_wt_mask_d_1_62;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_63 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_63 <= in_rt_wt_mask_d_1_63;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_64 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_64 <= in_rt_wt_mask_d_1_64;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_65 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_65 <= in_rt_wt_mask_d_1_65;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_66 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_66 <= in_rt_wt_mask_d_1_66;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_67 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_67 <= in_rt_wt_mask_d_1_67;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_68 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_68 <= in_rt_wt_mask_d_1_68;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_69 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_69 <= in_rt_wt_mask_d_1_69;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_70 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_70 <= in_rt_wt_mask_d_1_70;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_71 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_71 <= in_rt_wt_mask_d_1_71;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_72 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_72 <= in_rt_wt_mask_d_1_72;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_73 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_73 <= in_rt_wt_mask_d_1_73;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_74 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_74 <= in_rt_wt_mask_d_1_74;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_75 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_75 <= in_rt_wt_mask_d_1_75;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_76 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_76 <= in_rt_wt_mask_d_1_76;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_77 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_77 <= in_rt_wt_mask_d_1_77;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_78 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_78 <= in_rt_wt_mask_d_1_78;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_79 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_79 <= in_rt_wt_mask_d_1_79;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_80 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_80 <= in_rt_wt_mask_d_1_80;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_81 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_81 <= in_rt_wt_mask_d_1_81;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_82 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_82 <= in_rt_wt_mask_d_1_82;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_83 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_83 <= in_rt_wt_mask_d_1_83;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_84 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_84 <= in_rt_wt_mask_d_1_84;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_85 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_85 <= in_rt_wt_mask_d_1_85;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_86 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_86 <= in_rt_wt_mask_d_1_86;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_87 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_87 <= in_rt_wt_mask_d_1_87;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_88 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_88 <= in_rt_wt_mask_d_1_88;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_89 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_89 <= in_rt_wt_mask_d_1_89;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_90 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_90 <= in_rt_wt_mask_d_1_90;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_91 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_91 <= in_rt_wt_mask_d_1_91;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_92 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_92 <= in_rt_wt_mask_d_1_92;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_93 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_93 <= in_rt_wt_mask_d_1_93;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_94 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_94 <= in_rt_wt_mask_d_1_94;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_95 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_95 <= in_rt_wt_mask_d_1_95;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_96 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_96 <= in_rt_wt_mask_d_1_96;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_97 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_97 <= in_rt_wt_mask_d_1_97;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_98 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_98 <= in_rt_wt_mask_d_1_98;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_99 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_99 <= in_rt_wt_mask_d_1_99;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_100 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_100 <= in_rt_wt_mask_d_1_100;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_101 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_101 <= in_rt_wt_mask_d_1_101;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_102 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_102 <= in_rt_wt_mask_d_1_102;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_103 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_103 <= in_rt_wt_mask_d_1_103;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_104 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_104 <= in_rt_wt_mask_d_1_104;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_105 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_105 <= in_rt_wt_mask_d_1_105;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_106 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_106 <= in_rt_wt_mask_d_1_106;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_107 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_107 <= in_rt_wt_mask_d_1_107;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_108 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_108 <= in_rt_wt_mask_d_1_108;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_109 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_109 <= in_rt_wt_mask_d_1_109;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_110 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_110 <= in_rt_wt_mask_d_1_110;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_111 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_111 <= in_rt_wt_mask_d_1_111;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_112 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_112 <= in_rt_wt_mask_d_1_112;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_113 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_113 <= in_rt_wt_mask_d_1_113;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_114 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_114 <= in_rt_wt_mask_d_1_114;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_115 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_115 <= in_rt_wt_mask_d_1_115;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_116 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_116 <= in_rt_wt_mask_d_1_116;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_117 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_117 <= in_rt_wt_mask_d_1_117;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_118 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_118 <= in_rt_wt_mask_d_1_118;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_119 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_119 <= in_rt_wt_mask_d_1_119;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_120 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_120 <= in_rt_wt_mask_d_1_120;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_121 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_121 <= in_rt_wt_mask_d_1_121;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_122 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_122 <= in_rt_wt_mask_d_1_122;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_123 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_123 <= in_rt_wt_mask_d_1_123;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_124 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_124 <= in_rt_wt_mask_d_1_124;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_125 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_125 <= in_rt_wt_mask_d_1_125;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_126 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_126 <= in_rt_wt_mask_d_1_126;
      end
    end
    if (reset) begin
      in_rt_wt_mask_d_2_127 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_mask_d_2_127 <= in_rt_wt_mask_d_1_127;
      end
    end
    if (reset) begin
      in_rt_wt_pvld_d_1 <= 1'h0;
    end else begin
      in_rt_wt_pvld_d_1 <= io_sc2mac_wt_pvld;
    end
    if (reset) begin
      in_rt_wt_pvld_d_2 <= 1'h0;
    end else begin
      in_rt_wt_pvld_d_2 <= in_rt_wt_pvld_d_1;
    end
    if (reset) begin
      in_rt_wt_sel_d_1_0 <= 1'h0;
    end else begin
      if (_T_6929) begin
        in_rt_wt_sel_d_1_0 <= io_sc2mac_wt_sel_0;
      end
    end
    if (reset) begin
      in_rt_wt_sel_d_2_0 <= 1'h0;
    end else begin
      if (_T_6931) begin
        in_rt_wt_sel_d_2_0 <= in_rt_wt_sel_d_1_0;
      end
    end
  end
endmodule
module NV_NVDLA_CMAC_CORE_active(
  input        clock,
  input        reset,
  input  [7:0] io_in_dat_data_0,
  input  [7:0] io_in_dat_data_1,
  input  [7:0] io_in_dat_data_2,
  input  [7:0] io_in_dat_data_3,
  input  [7:0] io_in_dat_data_4,
  input  [7:0] io_in_dat_data_5,
  input  [7:0] io_in_dat_data_6,
  input  [7:0] io_in_dat_data_7,
  input  [7:0] io_in_dat_data_8,
  input  [7:0] io_in_dat_data_9,
  input  [7:0] io_in_dat_data_10,
  input  [7:0] io_in_dat_data_11,
  input  [7:0] io_in_dat_data_12,
  input  [7:0] io_in_dat_data_13,
  input  [7:0] io_in_dat_data_14,
  input  [7:0] io_in_dat_data_15,
  input  [7:0] io_in_dat_data_16,
  input  [7:0] io_in_dat_data_17,
  input  [7:0] io_in_dat_data_18,
  input  [7:0] io_in_dat_data_19,
  input  [7:0] io_in_dat_data_20,
  input  [7:0] io_in_dat_data_21,
  input  [7:0] io_in_dat_data_22,
  input  [7:0] io_in_dat_data_23,
  input  [7:0] io_in_dat_data_24,
  input  [7:0] io_in_dat_data_25,
  input  [7:0] io_in_dat_data_26,
  input  [7:0] io_in_dat_data_27,
  input  [7:0] io_in_dat_data_28,
  input  [7:0] io_in_dat_data_29,
  input  [7:0] io_in_dat_data_30,
  input  [7:0] io_in_dat_data_31,
  input  [7:0] io_in_dat_data_32,
  input  [7:0] io_in_dat_data_33,
  input  [7:0] io_in_dat_data_34,
  input  [7:0] io_in_dat_data_35,
  input  [7:0] io_in_dat_data_36,
  input  [7:0] io_in_dat_data_37,
  input  [7:0] io_in_dat_data_38,
  input  [7:0] io_in_dat_data_39,
  input  [7:0] io_in_dat_data_40,
  input  [7:0] io_in_dat_data_41,
  input  [7:0] io_in_dat_data_42,
  input  [7:0] io_in_dat_data_43,
  input  [7:0] io_in_dat_data_44,
  input  [7:0] io_in_dat_data_45,
  input  [7:0] io_in_dat_data_46,
  input  [7:0] io_in_dat_data_47,
  input  [7:0] io_in_dat_data_48,
  input  [7:0] io_in_dat_data_49,
  input  [7:0] io_in_dat_data_50,
  input  [7:0] io_in_dat_data_51,
  input  [7:0] io_in_dat_data_52,
  input  [7:0] io_in_dat_data_53,
  input  [7:0] io_in_dat_data_54,
  input  [7:0] io_in_dat_data_55,
  input  [7:0] io_in_dat_data_56,
  input  [7:0] io_in_dat_data_57,
  input  [7:0] io_in_dat_data_58,
  input  [7:0] io_in_dat_data_59,
  input  [7:0] io_in_dat_data_60,
  input  [7:0] io_in_dat_data_61,
  input  [7:0] io_in_dat_data_62,
  input  [7:0] io_in_dat_data_63,
  input  [7:0] io_in_dat_data_64,
  input  [7:0] io_in_dat_data_65,
  input  [7:0] io_in_dat_data_66,
  input  [7:0] io_in_dat_data_67,
  input  [7:0] io_in_dat_data_68,
  input  [7:0] io_in_dat_data_69,
  input  [7:0] io_in_dat_data_70,
  input  [7:0] io_in_dat_data_71,
  input  [7:0] io_in_dat_data_72,
  input  [7:0] io_in_dat_data_73,
  input  [7:0] io_in_dat_data_74,
  input  [7:0] io_in_dat_data_75,
  input  [7:0] io_in_dat_data_76,
  input  [7:0] io_in_dat_data_77,
  input  [7:0] io_in_dat_data_78,
  input  [7:0] io_in_dat_data_79,
  input  [7:0] io_in_dat_data_80,
  input  [7:0] io_in_dat_data_81,
  input  [7:0] io_in_dat_data_82,
  input  [7:0] io_in_dat_data_83,
  input  [7:0] io_in_dat_data_84,
  input  [7:0] io_in_dat_data_85,
  input  [7:0] io_in_dat_data_86,
  input  [7:0] io_in_dat_data_87,
  input  [7:0] io_in_dat_data_88,
  input  [7:0] io_in_dat_data_89,
  input  [7:0] io_in_dat_data_90,
  input  [7:0] io_in_dat_data_91,
  input  [7:0] io_in_dat_data_92,
  input  [7:0] io_in_dat_data_93,
  input  [7:0] io_in_dat_data_94,
  input  [7:0] io_in_dat_data_95,
  input  [7:0] io_in_dat_data_96,
  input  [7:0] io_in_dat_data_97,
  input  [7:0] io_in_dat_data_98,
  input  [7:0] io_in_dat_data_99,
  input  [7:0] io_in_dat_data_100,
  input  [7:0] io_in_dat_data_101,
  input  [7:0] io_in_dat_data_102,
  input  [7:0] io_in_dat_data_103,
  input  [7:0] io_in_dat_data_104,
  input  [7:0] io_in_dat_data_105,
  input  [7:0] io_in_dat_data_106,
  input  [7:0] io_in_dat_data_107,
  input  [7:0] io_in_dat_data_108,
  input  [7:0] io_in_dat_data_109,
  input  [7:0] io_in_dat_data_110,
  input  [7:0] io_in_dat_data_111,
  input  [7:0] io_in_dat_data_112,
  input  [7:0] io_in_dat_data_113,
  input  [7:0] io_in_dat_data_114,
  input  [7:0] io_in_dat_data_115,
  input  [7:0] io_in_dat_data_116,
  input  [7:0] io_in_dat_data_117,
  input  [7:0] io_in_dat_data_118,
  input  [7:0] io_in_dat_data_119,
  input  [7:0] io_in_dat_data_120,
  input  [7:0] io_in_dat_data_121,
  input  [7:0] io_in_dat_data_122,
  input  [7:0] io_in_dat_data_123,
  input  [7:0] io_in_dat_data_124,
  input  [7:0] io_in_dat_data_125,
  input  [7:0] io_in_dat_data_126,
  input  [7:0] io_in_dat_data_127,
  input        io_in_dat_mask_0,
  input        io_in_dat_mask_1,
  input        io_in_dat_mask_2,
  input        io_in_dat_mask_3,
  input        io_in_dat_mask_4,
  input        io_in_dat_mask_5,
  input        io_in_dat_mask_6,
  input        io_in_dat_mask_7,
  input        io_in_dat_mask_8,
  input        io_in_dat_mask_9,
  input        io_in_dat_mask_10,
  input        io_in_dat_mask_11,
  input        io_in_dat_mask_12,
  input        io_in_dat_mask_13,
  input        io_in_dat_mask_14,
  input        io_in_dat_mask_15,
  input        io_in_dat_mask_16,
  input        io_in_dat_mask_17,
  input        io_in_dat_mask_18,
  input        io_in_dat_mask_19,
  input        io_in_dat_mask_20,
  input        io_in_dat_mask_21,
  input        io_in_dat_mask_22,
  input        io_in_dat_mask_23,
  input        io_in_dat_mask_24,
  input        io_in_dat_mask_25,
  input        io_in_dat_mask_26,
  input        io_in_dat_mask_27,
  input        io_in_dat_mask_28,
  input        io_in_dat_mask_29,
  input        io_in_dat_mask_30,
  input        io_in_dat_mask_31,
  input        io_in_dat_mask_32,
  input        io_in_dat_mask_33,
  input        io_in_dat_mask_34,
  input        io_in_dat_mask_35,
  input        io_in_dat_mask_36,
  input        io_in_dat_mask_37,
  input        io_in_dat_mask_38,
  input        io_in_dat_mask_39,
  input        io_in_dat_mask_40,
  input        io_in_dat_mask_41,
  input        io_in_dat_mask_42,
  input        io_in_dat_mask_43,
  input        io_in_dat_mask_44,
  input        io_in_dat_mask_45,
  input        io_in_dat_mask_46,
  input        io_in_dat_mask_47,
  input        io_in_dat_mask_48,
  input        io_in_dat_mask_49,
  input        io_in_dat_mask_50,
  input        io_in_dat_mask_51,
  input        io_in_dat_mask_52,
  input        io_in_dat_mask_53,
  input        io_in_dat_mask_54,
  input        io_in_dat_mask_55,
  input        io_in_dat_mask_56,
  input        io_in_dat_mask_57,
  input        io_in_dat_mask_58,
  input        io_in_dat_mask_59,
  input        io_in_dat_mask_60,
  input        io_in_dat_mask_61,
  input        io_in_dat_mask_62,
  input        io_in_dat_mask_63,
  input        io_in_dat_mask_64,
  input        io_in_dat_mask_65,
  input        io_in_dat_mask_66,
  input        io_in_dat_mask_67,
  input        io_in_dat_mask_68,
  input        io_in_dat_mask_69,
  input        io_in_dat_mask_70,
  input        io_in_dat_mask_71,
  input        io_in_dat_mask_72,
  input        io_in_dat_mask_73,
  input        io_in_dat_mask_74,
  input        io_in_dat_mask_75,
  input        io_in_dat_mask_76,
  input        io_in_dat_mask_77,
  input        io_in_dat_mask_78,
  input        io_in_dat_mask_79,
  input        io_in_dat_mask_80,
  input        io_in_dat_mask_81,
  input        io_in_dat_mask_82,
  input        io_in_dat_mask_83,
  input        io_in_dat_mask_84,
  input        io_in_dat_mask_85,
  input        io_in_dat_mask_86,
  input        io_in_dat_mask_87,
  input        io_in_dat_mask_88,
  input        io_in_dat_mask_89,
  input        io_in_dat_mask_90,
  input        io_in_dat_mask_91,
  input        io_in_dat_mask_92,
  input        io_in_dat_mask_93,
  input        io_in_dat_mask_94,
  input        io_in_dat_mask_95,
  input        io_in_dat_mask_96,
  input        io_in_dat_mask_97,
  input        io_in_dat_mask_98,
  input        io_in_dat_mask_99,
  input        io_in_dat_mask_100,
  input        io_in_dat_mask_101,
  input        io_in_dat_mask_102,
  input        io_in_dat_mask_103,
  input        io_in_dat_mask_104,
  input        io_in_dat_mask_105,
  input        io_in_dat_mask_106,
  input        io_in_dat_mask_107,
  input        io_in_dat_mask_108,
  input        io_in_dat_mask_109,
  input        io_in_dat_mask_110,
  input        io_in_dat_mask_111,
  input        io_in_dat_mask_112,
  input        io_in_dat_mask_113,
  input        io_in_dat_mask_114,
  input        io_in_dat_mask_115,
  input        io_in_dat_mask_116,
  input        io_in_dat_mask_117,
  input        io_in_dat_mask_118,
  input        io_in_dat_mask_119,
  input        io_in_dat_mask_120,
  input        io_in_dat_mask_121,
  input        io_in_dat_mask_122,
  input        io_in_dat_mask_123,
  input        io_in_dat_mask_124,
  input        io_in_dat_mask_125,
  input        io_in_dat_mask_126,
  input        io_in_dat_mask_127,
  input        io_in_dat_pvld,
  input        io_in_dat_stripe_st,
  input        io_in_dat_stripe_end,
  input  [7:0] io_in_wt_data_0,
  input  [7:0] io_in_wt_data_1,
  input  [7:0] io_in_wt_data_2,
  input  [7:0] io_in_wt_data_3,
  input  [7:0] io_in_wt_data_4,
  input  [7:0] io_in_wt_data_5,
  input  [7:0] io_in_wt_data_6,
  input  [7:0] io_in_wt_data_7,
  input  [7:0] io_in_wt_data_8,
  input  [7:0] io_in_wt_data_9,
  input  [7:0] io_in_wt_data_10,
  input  [7:0] io_in_wt_data_11,
  input  [7:0] io_in_wt_data_12,
  input  [7:0] io_in_wt_data_13,
  input  [7:0] io_in_wt_data_14,
  input  [7:0] io_in_wt_data_15,
  input  [7:0] io_in_wt_data_16,
  input  [7:0] io_in_wt_data_17,
  input  [7:0] io_in_wt_data_18,
  input  [7:0] io_in_wt_data_19,
  input  [7:0] io_in_wt_data_20,
  input  [7:0] io_in_wt_data_21,
  input  [7:0] io_in_wt_data_22,
  input  [7:0] io_in_wt_data_23,
  input  [7:0] io_in_wt_data_24,
  input  [7:0] io_in_wt_data_25,
  input  [7:0] io_in_wt_data_26,
  input  [7:0] io_in_wt_data_27,
  input  [7:0] io_in_wt_data_28,
  input  [7:0] io_in_wt_data_29,
  input  [7:0] io_in_wt_data_30,
  input  [7:0] io_in_wt_data_31,
  input  [7:0] io_in_wt_data_32,
  input  [7:0] io_in_wt_data_33,
  input  [7:0] io_in_wt_data_34,
  input  [7:0] io_in_wt_data_35,
  input  [7:0] io_in_wt_data_36,
  input  [7:0] io_in_wt_data_37,
  input  [7:0] io_in_wt_data_38,
  input  [7:0] io_in_wt_data_39,
  input  [7:0] io_in_wt_data_40,
  input  [7:0] io_in_wt_data_41,
  input  [7:0] io_in_wt_data_42,
  input  [7:0] io_in_wt_data_43,
  input  [7:0] io_in_wt_data_44,
  input  [7:0] io_in_wt_data_45,
  input  [7:0] io_in_wt_data_46,
  input  [7:0] io_in_wt_data_47,
  input  [7:0] io_in_wt_data_48,
  input  [7:0] io_in_wt_data_49,
  input  [7:0] io_in_wt_data_50,
  input  [7:0] io_in_wt_data_51,
  input  [7:0] io_in_wt_data_52,
  input  [7:0] io_in_wt_data_53,
  input  [7:0] io_in_wt_data_54,
  input  [7:0] io_in_wt_data_55,
  input  [7:0] io_in_wt_data_56,
  input  [7:0] io_in_wt_data_57,
  input  [7:0] io_in_wt_data_58,
  input  [7:0] io_in_wt_data_59,
  input  [7:0] io_in_wt_data_60,
  input  [7:0] io_in_wt_data_61,
  input  [7:0] io_in_wt_data_62,
  input  [7:0] io_in_wt_data_63,
  input  [7:0] io_in_wt_data_64,
  input  [7:0] io_in_wt_data_65,
  input  [7:0] io_in_wt_data_66,
  input  [7:0] io_in_wt_data_67,
  input  [7:0] io_in_wt_data_68,
  input  [7:0] io_in_wt_data_69,
  input  [7:0] io_in_wt_data_70,
  input  [7:0] io_in_wt_data_71,
  input  [7:0] io_in_wt_data_72,
  input  [7:0] io_in_wt_data_73,
  input  [7:0] io_in_wt_data_74,
  input  [7:0] io_in_wt_data_75,
  input  [7:0] io_in_wt_data_76,
  input  [7:0] io_in_wt_data_77,
  input  [7:0] io_in_wt_data_78,
  input  [7:0] io_in_wt_data_79,
  input  [7:0] io_in_wt_data_80,
  input  [7:0] io_in_wt_data_81,
  input  [7:0] io_in_wt_data_82,
  input  [7:0] io_in_wt_data_83,
  input  [7:0] io_in_wt_data_84,
  input  [7:0] io_in_wt_data_85,
  input  [7:0] io_in_wt_data_86,
  input  [7:0] io_in_wt_data_87,
  input  [7:0] io_in_wt_data_88,
  input  [7:0] io_in_wt_data_89,
  input  [7:0] io_in_wt_data_90,
  input  [7:0] io_in_wt_data_91,
  input  [7:0] io_in_wt_data_92,
  input  [7:0] io_in_wt_data_93,
  input  [7:0] io_in_wt_data_94,
  input  [7:0] io_in_wt_data_95,
  input  [7:0] io_in_wt_data_96,
  input  [7:0] io_in_wt_data_97,
  input  [7:0] io_in_wt_data_98,
  input  [7:0] io_in_wt_data_99,
  input  [7:0] io_in_wt_data_100,
  input  [7:0] io_in_wt_data_101,
  input  [7:0] io_in_wt_data_102,
  input  [7:0] io_in_wt_data_103,
  input  [7:0] io_in_wt_data_104,
  input  [7:0] io_in_wt_data_105,
  input  [7:0] io_in_wt_data_106,
  input  [7:0] io_in_wt_data_107,
  input  [7:0] io_in_wt_data_108,
  input  [7:0] io_in_wt_data_109,
  input  [7:0] io_in_wt_data_110,
  input  [7:0] io_in_wt_data_111,
  input  [7:0] io_in_wt_data_112,
  input  [7:0] io_in_wt_data_113,
  input  [7:0] io_in_wt_data_114,
  input  [7:0] io_in_wt_data_115,
  input  [7:0] io_in_wt_data_116,
  input  [7:0] io_in_wt_data_117,
  input  [7:0] io_in_wt_data_118,
  input  [7:0] io_in_wt_data_119,
  input  [7:0] io_in_wt_data_120,
  input  [7:0] io_in_wt_data_121,
  input  [7:0] io_in_wt_data_122,
  input  [7:0] io_in_wt_data_123,
  input  [7:0] io_in_wt_data_124,
  input  [7:0] io_in_wt_data_125,
  input  [7:0] io_in_wt_data_126,
  input  [7:0] io_in_wt_data_127,
  input        io_in_wt_mask_0,
  input        io_in_wt_mask_1,
  input        io_in_wt_mask_2,
  input        io_in_wt_mask_3,
  input        io_in_wt_mask_4,
  input        io_in_wt_mask_5,
  input        io_in_wt_mask_6,
  input        io_in_wt_mask_7,
  input        io_in_wt_mask_8,
  input        io_in_wt_mask_9,
  input        io_in_wt_mask_10,
  input        io_in_wt_mask_11,
  input        io_in_wt_mask_12,
  input        io_in_wt_mask_13,
  input        io_in_wt_mask_14,
  input        io_in_wt_mask_15,
  input        io_in_wt_mask_16,
  input        io_in_wt_mask_17,
  input        io_in_wt_mask_18,
  input        io_in_wt_mask_19,
  input        io_in_wt_mask_20,
  input        io_in_wt_mask_21,
  input        io_in_wt_mask_22,
  input        io_in_wt_mask_23,
  input        io_in_wt_mask_24,
  input        io_in_wt_mask_25,
  input        io_in_wt_mask_26,
  input        io_in_wt_mask_27,
  input        io_in_wt_mask_28,
  input        io_in_wt_mask_29,
  input        io_in_wt_mask_30,
  input        io_in_wt_mask_31,
  input        io_in_wt_mask_32,
  input        io_in_wt_mask_33,
  input        io_in_wt_mask_34,
  input        io_in_wt_mask_35,
  input        io_in_wt_mask_36,
  input        io_in_wt_mask_37,
  input        io_in_wt_mask_38,
  input        io_in_wt_mask_39,
  input        io_in_wt_mask_40,
  input        io_in_wt_mask_41,
  input        io_in_wt_mask_42,
  input        io_in_wt_mask_43,
  input        io_in_wt_mask_44,
  input        io_in_wt_mask_45,
  input        io_in_wt_mask_46,
  input        io_in_wt_mask_47,
  input        io_in_wt_mask_48,
  input        io_in_wt_mask_49,
  input        io_in_wt_mask_50,
  input        io_in_wt_mask_51,
  input        io_in_wt_mask_52,
  input        io_in_wt_mask_53,
  input        io_in_wt_mask_54,
  input        io_in_wt_mask_55,
  input        io_in_wt_mask_56,
  input        io_in_wt_mask_57,
  input        io_in_wt_mask_58,
  input        io_in_wt_mask_59,
  input        io_in_wt_mask_60,
  input        io_in_wt_mask_61,
  input        io_in_wt_mask_62,
  input        io_in_wt_mask_63,
  input        io_in_wt_mask_64,
  input        io_in_wt_mask_65,
  input        io_in_wt_mask_66,
  input        io_in_wt_mask_67,
  input        io_in_wt_mask_68,
  input        io_in_wt_mask_69,
  input        io_in_wt_mask_70,
  input        io_in_wt_mask_71,
  input        io_in_wt_mask_72,
  input        io_in_wt_mask_73,
  input        io_in_wt_mask_74,
  input        io_in_wt_mask_75,
  input        io_in_wt_mask_76,
  input        io_in_wt_mask_77,
  input        io_in_wt_mask_78,
  input        io_in_wt_mask_79,
  input        io_in_wt_mask_80,
  input        io_in_wt_mask_81,
  input        io_in_wt_mask_82,
  input        io_in_wt_mask_83,
  input        io_in_wt_mask_84,
  input        io_in_wt_mask_85,
  input        io_in_wt_mask_86,
  input        io_in_wt_mask_87,
  input        io_in_wt_mask_88,
  input        io_in_wt_mask_89,
  input        io_in_wt_mask_90,
  input        io_in_wt_mask_91,
  input        io_in_wt_mask_92,
  input        io_in_wt_mask_93,
  input        io_in_wt_mask_94,
  input        io_in_wt_mask_95,
  input        io_in_wt_mask_96,
  input        io_in_wt_mask_97,
  input        io_in_wt_mask_98,
  input        io_in_wt_mask_99,
  input        io_in_wt_mask_100,
  input        io_in_wt_mask_101,
  input        io_in_wt_mask_102,
  input        io_in_wt_mask_103,
  input        io_in_wt_mask_104,
  input        io_in_wt_mask_105,
  input        io_in_wt_mask_106,
  input        io_in_wt_mask_107,
  input        io_in_wt_mask_108,
  input        io_in_wt_mask_109,
  input        io_in_wt_mask_110,
  input        io_in_wt_mask_111,
  input        io_in_wt_mask_112,
  input        io_in_wt_mask_113,
  input        io_in_wt_mask_114,
  input        io_in_wt_mask_115,
  input        io_in_wt_mask_116,
  input        io_in_wt_mask_117,
  input        io_in_wt_mask_118,
  input        io_in_wt_mask_119,
  input        io_in_wt_mask_120,
  input        io_in_wt_mask_121,
  input        io_in_wt_mask_122,
  input        io_in_wt_mask_123,
  input        io_in_wt_mask_124,
  input        io_in_wt_mask_125,
  input        io_in_wt_mask_126,
  input        io_in_wt_mask_127,
  input        io_in_wt_pvld,
  input        io_in_wt_sel_0,
  output [7:0] io_dat_actv_data_0_0,
  output [7:0] io_dat_actv_data_0_1,
  output [7:0] io_dat_actv_data_0_2,
  output [7:0] io_dat_actv_data_0_3,
  output [7:0] io_dat_actv_data_0_4,
  output [7:0] io_dat_actv_data_0_5,
  output [7:0] io_dat_actv_data_0_6,
  output [7:0] io_dat_actv_data_0_7,
  output [7:0] io_dat_actv_data_0_8,
  output [7:0] io_dat_actv_data_0_9,
  output [7:0] io_dat_actv_data_0_10,
  output [7:0] io_dat_actv_data_0_11,
  output [7:0] io_dat_actv_data_0_12,
  output [7:0] io_dat_actv_data_0_13,
  output [7:0] io_dat_actv_data_0_14,
  output [7:0] io_dat_actv_data_0_15,
  output [7:0] io_dat_actv_data_0_16,
  output [7:0] io_dat_actv_data_0_17,
  output [7:0] io_dat_actv_data_0_18,
  output [7:0] io_dat_actv_data_0_19,
  output [7:0] io_dat_actv_data_0_20,
  output [7:0] io_dat_actv_data_0_21,
  output [7:0] io_dat_actv_data_0_22,
  output [7:0] io_dat_actv_data_0_23,
  output [7:0] io_dat_actv_data_0_24,
  output [7:0] io_dat_actv_data_0_25,
  output [7:0] io_dat_actv_data_0_26,
  output [7:0] io_dat_actv_data_0_27,
  output [7:0] io_dat_actv_data_0_28,
  output [7:0] io_dat_actv_data_0_29,
  output [7:0] io_dat_actv_data_0_30,
  output [7:0] io_dat_actv_data_0_31,
  output [7:0] io_dat_actv_data_0_32,
  output [7:0] io_dat_actv_data_0_33,
  output [7:0] io_dat_actv_data_0_34,
  output [7:0] io_dat_actv_data_0_35,
  output [7:0] io_dat_actv_data_0_36,
  output [7:0] io_dat_actv_data_0_37,
  output [7:0] io_dat_actv_data_0_38,
  output [7:0] io_dat_actv_data_0_39,
  output [7:0] io_dat_actv_data_0_40,
  output [7:0] io_dat_actv_data_0_41,
  output [7:0] io_dat_actv_data_0_42,
  output [7:0] io_dat_actv_data_0_43,
  output [7:0] io_dat_actv_data_0_44,
  output [7:0] io_dat_actv_data_0_45,
  output [7:0] io_dat_actv_data_0_46,
  output [7:0] io_dat_actv_data_0_47,
  output [7:0] io_dat_actv_data_0_48,
  output [7:0] io_dat_actv_data_0_49,
  output [7:0] io_dat_actv_data_0_50,
  output [7:0] io_dat_actv_data_0_51,
  output [7:0] io_dat_actv_data_0_52,
  output [7:0] io_dat_actv_data_0_53,
  output [7:0] io_dat_actv_data_0_54,
  output [7:0] io_dat_actv_data_0_55,
  output [7:0] io_dat_actv_data_0_56,
  output [7:0] io_dat_actv_data_0_57,
  output [7:0] io_dat_actv_data_0_58,
  output [7:0] io_dat_actv_data_0_59,
  output [7:0] io_dat_actv_data_0_60,
  output [7:0] io_dat_actv_data_0_61,
  output [7:0] io_dat_actv_data_0_62,
  output [7:0] io_dat_actv_data_0_63,
  output [7:0] io_dat_actv_data_0_64,
  output [7:0] io_dat_actv_data_0_65,
  output [7:0] io_dat_actv_data_0_66,
  output [7:0] io_dat_actv_data_0_67,
  output [7:0] io_dat_actv_data_0_68,
  output [7:0] io_dat_actv_data_0_69,
  output [7:0] io_dat_actv_data_0_70,
  output [7:0] io_dat_actv_data_0_71,
  output [7:0] io_dat_actv_data_0_72,
  output [7:0] io_dat_actv_data_0_73,
  output [7:0] io_dat_actv_data_0_74,
  output [7:0] io_dat_actv_data_0_75,
  output [7:0] io_dat_actv_data_0_76,
  output [7:0] io_dat_actv_data_0_77,
  output [7:0] io_dat_actv_data_0_78,
  output [7:0] io_dat_actv_data_0_79,
  output [7:0] io_dat_actv_data_0_80,
  output [7:0] io_dat_actv_data_0_81,
  output [7:0] io_dat_actv_data_0_82,
  output [7:0] io_dat_actv_data_0_83,
  output [7:0] io_dat_actv_data_0_84,
  output [7:0] io_dat_actv_data_0_85,
  output [7:0] io_dat_actv_data_0_86,
  output [7:0] io_dat_actv_data_0_87,
  output [7:0] io_dat_actv_data_0_88,
  output [7:0] io_dat_actv_data_0_89,
  output [7:0] io_dat_actv_data_0_90,
  output [7:0] io_dat_actv_data_0_91,
  output [7:0] io_dat_actv_data_0_92,
  output [7:0] io_dat_actv_data_0_93,
  output [7:0] io_dat_actv_data_0_94,
  output [7:0] io_dat_actv_data_0_95,
  output [7:0] io_dat_actv_data_0_96,
  output [7:0] io_dat_actv_data_0_97,
  output [7:0] io_dat_actv_data_0_98,
  output [7:0] io_dat_actv_data_0_99,
  output [7:0] io_dat_actv_data_0_100,
  output [7:0] io_dat_actv_data_0_101,
  output [7:0] io_dat_actv_data_0_102,
  output [7:0] io_dat_actv_data_0_103,
  output [7:0] io_dat_actv_data_0_104,
  output [7:0] io_dat_actv_data_0_105,
  output [7:0] io_dat_actv_data_0_106,
  output [7:0] io_dat_actv_data_0_107,
  output [7:0] io_dat_actv_data_0_108,
  output [7:0] io_dat_actv_data_0_109,
  output [7:0] io_dat_actv_data_0_110,
  output [7:0] io_dat_actv_data_0_111,
  output [7:0] io_dat_actv_data_0_112,
  output [7:0] io_dat_actv_data_0_113,
  output [7:0] io_dat_actv_data_0_114,
  output [7:0] io_dat_actv_data_0_115,
  output [7:0] io_dat_actv_data_0_116,
  output [7:0] io_dat_actv_data_0_117,
  output [7:0] io_dat_actv_data_0_118,
  output [7:0] io_dat_actv_data_0_119,
  output [7:0] io_dat_actv_data_0_120,
  output [7:0] io_dat_actv_data_0_121,
  output [7:0] io_dat_actv_data_0_122,
  output [7:0] io_dat_actv_data_0_123,
  output [7:0] io_dat_actv_data_0_124,
  output [7:0] io_dat_actv_data_0_125,
  output [7:0] io_dat_actv_data_0_126,
  output [7:0] io_dat_actv_data_0_127,
  output       io_dat_actv_nz_0_0,
  output       io_dat_actv_nz_0_1,
  output       io_dat_actv_nz_0_2,
  output       io_dat_actv_nz_0_3,
  output       io_dat_actv_nz_0_4,
  output       io_dat_actv_nz_0_5,
  output       io_dat_actv_nz_0_6,
  output       io_dat_actv_nz_0_7,
  output       io_dat_actv_nz_0_8,
  output       io_dat_actv_nz_0_9,
  output       io_dat_actv_nz_0_10,
  output       io_dat_actv_nz_0_11,
  output       io_dat_actv_nz_0_12,
  output       io_dat_actv_nz_0_13,
  output       io_dat_actv_nz_0_14,
  output       io_dat_actv_nz_0_15,
  output       io_dat_actv_nz_0_16,
  output       io_dat_actv_nz_0_17,
  output       io_dat_actv_nz_0_18,
  output       io_dat_actv_nz_0_19,
  output       io_dat_actv_nz_0_20,
  output       io_dat_actv_nz_0_21,
  output       io_dat_actv_nz_0_22,
  output       io_dat_actv_nz_0_23,
  output       io_dat_actv_nz_0_24,
  output       io_dat_actv_nz_0_25,
  output       io_dat_actv_nz_0_26,
  output       io_dat_actv_nz_0_27,
  output       io_dat_actv_nz_0_28,
  output       io_dat_actv_nz_0_29,
  output       io_dat_actv_nz_0_30,
  output       io_dat_actv_nz_0_31,
  output       io_dat_actv_nz_0_32,
  output       io_dat_actv_nz_0_33,
  output       io_dat_actv_nz_0_34,
  output       io_dat_actv_nz_0_35,
  output       io_dat_actv_nz_0_36,
  output       io_dat_actv_nz_0_37,
  output       io_dat_actv_nz_0_38,
  output       io_dat_actv_nz_0_39,
  output       io_dat_actv_nz_0_40,
  output       io_dat_actv_nz_0_41,
  output       io_dat_actv_nz_0_42,
  output       io_dat_actv_nz_0_43,
  output       io_dat_actv_nz_0_44,
  output       io_dat_actv_nz_0_45,
  output       io_dat_actv_nz_0_46,
  output       io_dat_actv_nz_0_47,
  output       io_dat_actv_nz_0_48,
  output       io_dat_actv_nz_0_49,
  output       io_dat_actv_nz_0_50,
  output       io_dat_actv_nz_0_51,
  output       io_dat_actv_nz_0_52,
  output       io_dat_actv_nz_0_53,
  output       io_dat_actv_nz_0_54,
  output       io_dat_actv_nz_0_55,
  output       io_dat_actv_nz_0_56,
  output       io_dat_actv_nz_0_57,
  output       io_dat_actv_nz_0_58,
  output       io_dat_actv_nz_0_59,
  output       io_dat_actv_nz_0_60,
  output       io_dat_actv_nz_0_61,
  output       io_dat_actv_nz_0_62,
  output       io_dat_actv_nz_0_63,
  output       io_dat_actv_nz_0_64,
  output       io_dat_actv_nz_0_65,
  output       io_dat_actv_nz_0_66,
  output       io_dat_actv_nz_0_67,
  output       io_dat_actv_nz_0_68,
  output       io_dat_actv_nz_0_69,
  output       io_dat_actv_nz_0_70,
  output       io_dat_actv_nz_0_71,
  output       io_dat_actv_nz_0_72,
  output       io_dat_actv_nz_0_73,
  output       io_dat_actv_nz_0_74,
  output       io_dat_actv_nz_0_75,
  output       io_dat_actv_nz_0_76,
  output       io_dat_actv_nz_0_77,
  output       io_dat_actv_nz_0_78,
  output       io_dat_actv_nz_0_79,
  output       io_dat_actv_nz_0_80,
  output       io_dat_actv_nz_0_81,
  output       io_dat_actv_nz_0_82,
  output       io_dat_actv_nz_0_83,
  output       io_dat_actv_nz_0_84,
  output       io_dat_actv_nz_0_85,
  output       io_dat_actv_nz_0_86,
  output       io_dat_actv_nz_0_87,
  output       io_dat_actv_nz_0_88,
  output       io_dat_actv_nz_0_89,
  output       io_dat_actv_nz_0_90,
  output       io_dat_actv_nz_0_91,
  output       io_dat_actv_nz_0_92,
  output       io_dat_actv_nz_0_93,
  output       io_dat_actv_nz_0_94,
  output       io_dat_actv_nz_0_95,
  output       io_dat_actv_nz_0_96,
  output       io_dat_actv_nz_0_97,
  output       io_dat_actv_nz_0_98,
  output       io_dat_actv_nz_0_99,
  output       io_dat_actv_nz_0_100,
  output       io_dat_actv_nz_0_101,
  output       io_dat_actv_nz_0_102,
  output       io_dat_actv_nz_0_103,
  output       io_dat_actv_nz_0_104,
  output       io_dat_actv_nz_0_105,
  output       io_dat_actv_nz_0_106,
  output       io_dat_actv_nz_0_107,
  output       io_dat_actv_nz_0_108,
  output       io_dat_actv_nz_0_109,
  output       io_dat_actv_nz_0_110,
  output       io_dat_actv_nz_0_111,
  output       io_dat_actv_nz_0_112,
  output       io_dat_actv_nz_0_113,
  output       io_dat_actv_nz_0_114,
  output       io_dat_actv_nz_0_115,
  output       io_dat_actv_nz_0_116,
  output       io_dat_actv_nz_0_117,
  output       io_dat_actv_nz_0_118,
  output       io_dat_actv_nz_0_119,
  output       io_dat_actv_nz_0_120,
  output       io_dat_actv_nz_0_121,
  output       io_dat_actv_nz_0_122,
  output       io_dat_actv_nz_0_123,
  output       io_dat_actv_nz_0_124,
  output       io_dat_actv_nz_0_125,
  output       io_dat_actv_nz_0_126,
  output       io_dat_actv_nz_0_127,
  output       io_dat_actv_pvld_0_0,
  output       io_dat_actv_pvld_0_1,
  output       io_dat_actv_pvld_0_2,
  output       io_dat_actv_pvld_0_3,
  output       io_dat_actv_pvld_0_4,
  output       io_dat_actv_pvld_0_5,
  output       io_dat_actv_pvld_0_6,
  output       io_dat_actv_pvld_0_7,
  output       io_dat_actv_pvld_0_8,
  output       io_dat_actv_pvld_0_9,
  output       io_dat_actv_pvld_0_10,
  output       io_dat_actv_pvld_0_11,
  output       io_dat_actv_pvld_0_12,
  output       io_dat_actv_pvld_0_13,
  output       io_dat_actv_pvld_0_14,
  output       io_dat_actv_pvld_0_15,
  output       io_dat_actv_pvld_0_16,
  output       io_dat_actv_pvld_0_17,
  output       io_dat_actv_pvld_0_18,
  output       io_dat_actv_pvld_0_19,
  output       io_dat_actv_pvld_0_20,
  output       io_dat_actv_pvld_0_21,
  output       io_dat_actv_pvld_0_22,
  output       io_dat_actv_pvld_0_23,
  output       io_dat_actv_pvld_0_24,
  output       io_dat_actv_pvld_0_25,
  output       io_dat_actv_pvld_0_26,
  output       io_dat_actv_pvld_0_27,
  output       io_dat_actv_pvld_0_28,
  output       io_dat_actv_pvld_0_29,
  output       io_dat_actv_pvld_0_30,
  output       io_dat_actv_pvld_0_31,
  output       io_dat_actv_pvld_0_32,
  output       io_dat_actv_pvld_0_33,
  output       io_dat_actv_pvld_0_34,
  output       io_dat_actv_pvld_0_35,
  output       io_dat_actv_pvld_0_36,
  output       io_dat_actv_pvld_0_37,
  output       io_dat_actv_pvld_0_38,
  output       io_dat_actv_pvld_0_39,
  output       io_dat_actv_pvld_0_40,
  output       io_dat_actv_pvld_0_41,
  output       io_dat_actv_pvld_0_42,
  output       io_dat_actv_pvld_0_43,
  output       io_dat_actv_pvld_0_44,
  output       io_dat_actv_pvld_0_45,
  output       io_dat_actv_pvld_0_46,
  output       io_dat_actv_pvld_0_47,
  output       io_dat_actv_pvld_0_48,
  output       io_dat_actv_pvld_0_49,
  output       io_dat_actv_pvld_0_50,
  output       io_dat_actv_pvld_0_51,
  output       io_dat_actv_pvld_0_52,
  output       io_dat_actv_pvld_0_53,
  output       io_dat_actv_pvld_0_54,
  output       io_dat_actv_pvld_0_55,
  output       io_dat_actv_pvld_0_56,
  output       io_dat_actv_pvld_0_57,
  output       io_dat_actv_pvld_0_58,
  output       io_dat_actv_pvld_0_59,
  output       io_dat_actv_pvld_0_60,
  output       io_dat_actv_pvld_0_61,
  output       io_dat_actv_pvld_0_62,
  output       io_dat_actv_pvld_0_63,
  output       io_dat_actv_pvld_0_64,
  output       io_dat_actv_pvld_0_65,
  output       io_dat_actv_pvld_0_66,
  output       io_dat_actv_pvld_0_67,
  output       io_dat_actv_pvld_0_68,
  output       io_dat_actv_pvld_0_69,
  output       io_dat_actv_pvld_0_70,
  output       io_dat_actv_pvld_0_71,
  output       io_dat_actv_pvld_0_72,
  output       io_dat_actv_pvld_0_73,
  output       io_dat_actv_pvld_0_74,
  output       io_dat_actv_pvld_0_75,
  output       io_dat_actv_pvld_0_76,
  output       io_dat_actv_pvld_0_77,
  output       io_dat_actv_pvld_0_78,
  output       io_dat_actv_pvld_0_79,
  output       io_dat_actv_pvld_0_80,
  output       io_dat_actv_pvld_0_81,
  output       io_dat_actv_pvld_0_82,
  output       io_dat_actv_pvld_0_83,
  output       io_dat_actv_pvld_0_84,
  output       io_dat_actv_pvld_0_85,
  output       io_dat_actv_pvld_0_86,
  output       io_dat_actv_pvld_0_87,
  output       io_dat_actv_pvld_0_88,
  output       io_dat_actv_pvld_0_89,
  output       io_dat_actv_pvld_0_90,
  output       io_dat_actv_pvld_0_91,
  output       io_dat_actv_pvld_0_92,
  output       io_dat_actv_pvld_0_93,
  output       io_dat_actv_pvld_0_94,
  output       io_dat_actv_pvld_0_95,
  output       io_dat_actv_pvld_0_96,
  output       io_dat_actv_pvld_0_97,
  output       io_dat_actv_pvld_0_98,
  output       io_dat_actv_pvld_0_99,
  output       io_dat_actv_pvld_0_100,
  output       io_dat_actv_pvld_0_101,
  output       io_dat_actv_pvld_0_102,
  output       io_dat_actv_pvld_0_103,
  output       io_dat_actv_pvld_0_104,
  output       io_dat_actv_pvld_0_105,
  output       io_dat_actv_pvld_0_106,
  output       io_dat_actv_pvld_0_107,
  output       io_dat_actv_pvld_0_108,
  output       io_dat_actv_pvld_0_109,
  output       io_dat_actv_pvld_0_110,
  output       io_dat_actv_pvld_0_111,
  output       io_dat_actv_pvld_0_112,
  output       io_dat_actv_pvld_0_113,
  output       io_dat_actv_pvld_0_114,
  output       io_dat_actv_pvld_0_115,
  output       io_dat_actv_pvld_0_116,
  output       io_dat_actv_pvld_0_117,
  output       io_dat_actv_pvld_0_118,
  output       io_dat_actv_pvld_0_119,
  output       io_dat_actv_pvld_0_120,
  output       io_dat_actv_pvld_0_121,
  output       io_dat_actv_pvld_0_122,
  output       io_dat_actv_pvld_0_123,
  output       io_dat_actv_pvld_0_124,
  output       io_dat_actv_pvld_0_125,
  output       io_dat_actv_pvld_0_126,
  output       io_dat_actv_pvld_0_127,
  output [7:0] io_wt_actv_data_0_0,
  output [7:0] io_wt_actv_data_0_1,
  output [7:0] io_wt_actv_data_0_2,
  output [7:0] io_wt_actv_data_0_3,
  output [7:0] io_wt_actv_data_0_4,
  output [7:0] io_wt_actv_data_0_5,
  output [7:0] io_wt_actv_data_0_6,
  output [7:0] io_wt_actv_data_0_7,
  output [7:0] io_wt_actv_data_0_8,
  output [7:0] io_wt_actv_data_0_9,
  output [7:0] io_wt_actv_data_0_10,
  output [7:0] io_wt_actv_data_0_11,
  output [7:0] io_wt_actv_data_0_12,
  output [7:0] io_wt_actv_data_0_13,
  output [7:0] io_wt_actv_data_0_14,
  output [7:0] io_wt_actv_data_0_15,
  output [7:0] io_wt_actv_data_0_16,
  output [7:0] io_wt_actv_data_0_17,
  output [7:0] io_wt_actv_data_0_18,
  output [7:0] io_wt_actv_data_0_19,
  output [7:0] io_wt_actv_data_0_20,
  output [7:0] io_wt_actv_data_0_21,
  output [7:0] io_wt_actv_data_0_22,
  output [7:0] io_wt_actv_data_0_23,
  output [7:0] io_wt_actv_data_0_24,
  output [7:0] io_wt_actv_data_0_25,
  output [7:0] io_wt_actv_data_0_26,
  output [7:0] io_wt_actv_data_0_27,
  output [7:0] io_wt_actv_data_0_28,
  output [7:0] io_wt_actv_data_0_29,
  output [7:0] io_wt_actv_data_0_30,
  output [7:0] io_wt_actv_data_0_31,
  output [7:0] io_wt_actv_data_0_32,
  output [7:0] io_wt_actv_data_0_33,
  output [7:0] io_wt_actv_data_0_34,
  output [7:0] io_wt_actv_data_0_35,
  output [7:0] io_wt_actv_data_0_36,
  output [7:0] io_wt_actv_data_0_37,
  output [7:0] io_wt_actv_data_0_38,
  output [7:0] io_wt_actv_data_0_39,
  output [7:0] io_wt_actv_data_0_40,
  output [7:0] io_wt_actv_data_0_41,
  output [7:0] io_wt_actv_data_0_42,
  output [7:0] io_wt_actv_data_0_43,
  output [7:0] io_wt_actv_data_0_44,
  output [7:0] io_wt_actv_data_0_45,
  output [7:0] io_wt_actv_data_0_46,
  output [7:0] io_wt_actv_data_0_47,
  output [7:0] io_wt_actv_data_0_48,
  output [7:0] io_wt_actv_data_0_49,
  output [7:0] io_wt_actv_data_0_50,
  output [7:0] io_wt_actv_data_0_51,
  output [7:0] io_wt_actv_data_0_52,
  output [7:0] io_wt_actv_data_0_53,
  output [7:0] io_wt_actv_data_0_54,
  output [7:0] io_wt_actv_data_0_55,
  output [7:0] io_wt_actv_data_0_56,
  output [7:0] io_wt_actv_data_0_57,
  output [7:0] io_wt_actv_data_0_58,
  output [7:0] io_wt_actv_data_0_59,
  output [7:0] io_wt_actv_data_0_60,
  output [7:0] io_wt_actv_data_0_61,
  output [7:0] io_wt_actv_data_0_62,
  output [7:0] io_wt_actv_data_0_63,
  output [7:0] io_wt_actv_data_0_64,
  output [7:0] io_wt_actv_data_0_65,
  output [7:0] io_wt_actv_data_0_66,
  output [7:0] io_wt_actv_data_0_67,
  output [7:0] io_wt_actv_data_0_68,
  output [7:0] io_wt_actv_data_0_69,
  output [7:0] io_wt_actv_data_0_70,
  output [7:0] io_wt_actv_data_0_71,
  output [7:0] io_wt_actv_data_0_72,
  output [7:0] io_wt_actv_data_0_73,
  output [7:0] io_wt_actv_data_0_74,
  output [7:0] io_wt_actv_data_0_75,
  output [7:0] io_wt_actv_data_0_76,
  output [7:0] io_wt_actv_data_0_77,
  output [7:0] io_wt_actv_data_0_78,
  output [7:0] io_wt_actv_data_0_79,
  output [7:0] io_wt_actv_data_0_80,
  output [7:0] io_wt_actv_data_0_81,
  output [7:0] io_wt_actv_data_0_82,
  output [7:0] io_wt_actv_data_0_83,
  output [7:0] io_wt_actv_data_0_84,
  output [7:0] io_wt_actv_data_0_85,
  output [7:0] io_wt_actv_data_0_86,
  output [7:0] io_wt_actv_data_0_87,
  output [7:0] io_wt_actv_data_0_88,
  output [7:0] io_wt_actv_data_0_89,
  output [7:0] io_wt_actv_data_0_90,
  output [7:0] io_wt_actv_data_0_91,
  output [7:0] io_wt_actv_data_0_92,
  output [7:0] io_wt_actv_data_0_93,
  output [7:0] io_wt_actv_data_0_94,
  output [7:0] io_wt_actv_data_0_95,
  output [7:0] io_wt_actv_data_0_96,
  output [7:0] io_wt_actv_data_0_97,
  output [7:0] io_wt_actv_data_0_98,
  output [7:0] io_wt_actv_data_0_99,
  output [7:0] io_wt_actv_data_0_100,
  output [7:0] io_wt_actv_data_0_101,
  output [7:0] io_wt_actv_data_0_102,
  output [7:0] io_wt_actv_data_0_103,
  output [7:0] io_wt_actv_data_0_104,
  output [7:0] io_wt_actv_data_0_105,
  output [7:0] io_wt_actv_data_0_106,
  output [7:0] io_wt_actv_data_0_107,
  output [7:0] io_wt_actv_data_0_108,
  output [7:0] io_wt_actv_data_0_109,
  output [7:0] io_wt_actv_data_0_110,
  output [7:0] io_wt_actv_data_0_111,
  output [7:0] io_wt_actv_data_0_112,
  output [7:0] io_wt_actv_data_0_113,
  output [7:0] io_wt_actv_data_0_114,
  output [7:0] io_wt_actv_data_0_115,
  output [7:0] io_wt_actv_data_0_116,
  output [7:0] io_wt_actv_data_0_117,
  output [7:0] io_wt_actv_data_0_118,
  output [7:0] io_wt_actv_data_0_119,
  output [7:0] io_wt_actv_data_0_120,
  output [7:0] io_wt_actv_data_0_121,
  output [7:0] io_wt_actv_data_0_122,
  output [7:0] io_wt_actv_data_0_123,
  output [7:0] io_wt_actv_data_0_124,
  output [7:0] io_wt_actv_data_0_125,
  output [7:0] io_wt_actv_data_0_126,
  output [7:0] io_wt_actv_data_0_127,
  output       io_wt_actv_nz_0_0,
  output       io_wt_actv_nz_0_1,
  output       io_wt_actv_nz_0_2,
  output       io_wt_actv_nz_0_3,
  output       io_wt_actv_nz_0_4,
  output       io_wt_actv_nz_0_5,
  output       io_wt_actv_nz_0_6,
  output       io_wt_actv_nz_0_7,
  output       io_wt_actv_nz_0_8,
  output       io_wt_actv_nz_0_9,
  output       io_wt_actv_nz_0_10,
  output       io_wt_actv_nz_0_11,
  output       io_wt_actv_nz_0_12,
  output       io_wt_actv_nz_0_13,
  output       io_wt_actv_nz_0_14,
  output       io_wt_actv_nz_0_15,
  output       io_wt_actv_nz_0_16,
  output       io_wt_actv_nz_0_17,
  output       io_wt_actv_nz_0_18,
  output       io_wt_actv_nz_0_19,
  output       io_wt_actv_nz_0_20,
  output       io_wt_actv_nz_0_21,
  output       io_wt_actv_nz_0_22,
  output       io_wt_actv_nz_0_23,
  output       io_wt_actv_nz_0_24,
  output       io_wt_actv_nz_0_25,
  output       io_wt_actv_nz_0_26,
  output       io_wt_actv_nz_0_27,
  output       io_wt_actv_nz_0_28,
  output       io_wt_actv_nz_0_29,
  output       io_wt_actv_nz_0_30,
  output       io_wt_actv_nz_0_31,
  output       io_wt_actv_nz_0_32,
  output       io_wt_actv_nz_0_33,
  output       io_wt_actv_nz_0_34,
  output       io_wt_actv_nz_0_35,
  output       io_wt_actv_nz_0_36,
  output       io_wt_actv_nz_0_37,
  output       io_wt_actv_nz_0_38,
  output       io_wt_actv_nz_0_39,
  output       io_wt_actv_nz_0_40,
  output       io_wt_actv_nz_0_41,
  output       io_wt_actv_nz_0_42,
  output       io_wt_actv_nz_0_43,
  output       io_wt_actv_nz_0_44,
  output       io_wt_actv_nz_0_45,
  output       io_wt_actv_nz_0_46,
  output       io_wt_actv_nz_0_47,
  output       io_wt_actv_nz_0_48,
  output       io_wt_actv_nz_0_49,
  output       io_wt_actv_nz_0_50,
  output       io_wt_actv_nz_0_51,
  output       io_wt_actv_nz_0_52,
  output       io_wt_actv_nz_0_53,
  output       io_wt_actv_nz_0_54,
  output       io_wt_actv_nz_0_55,
  output       io_wt_actv_nz_0_56,
  output       io_wt_actv_nz_0_57,
  output       io_wt_actv_nz_0_58,
  output       io_wt_actv_nz_0_59,
  output       io_wt_actv_nz_0_60,
  output       io_wt_actv_nz_0_61,
  output       io_wt_actv_nz_0_62,
  output       io_wt_actv_nz_0_63,
  output       io_wt_actv_nz_0_64,
  output       io_wt_actv_nz_0_65,
  output       io_wt_actv_nz_0_66,
  output       io_wt_actv_nz_0_67,
  output       io_wt_actv_nz_0_68,
  output       io_wt_actv_nz_0_69,
  output       io_wt_actv_nz_0_70,
  output       io_wt_actv_nz_0_71,
  output       io_wt_actv_nz_0_72,
  output       io_wt_actv_nz_0_73,
  output       io_wt_actv_nz_0_74,
  output       io_wt_actv_nz_0_75,
  output       io_wt_actv_nz_0_76,
  output       io_wt_actv_nz_0_77,
  output       io_wt_actv_nz_0_78,
  output       io_wt_actv_nz_0_79,
  output       io_wt_actv_nz_0_80,
  output       io_wt_actv_nz_0_81,
  output       io_wt_actv_nz_0_82,
  output       io_wt_actv_nz_0_83,
  output       io_wt_actv_nz_0_84,
  output       io_wt_actv_nz_0_85,
  output       io_wt_actv_nz_0_86,
  output       io_wt_actv_nz_0_87,
  output       io_wt_actv_nz_0_88,
  output       io_wt_actv_nz_0_89,
  output       io_wt_actv_nz_0_90,
  output       io_wt_actv_nz_0_91,
  output       io_wt_actv_nz_0_92,
  output       io_wt_actv_nz_0_93,
  output       io_wt_actv_nz_0_94,
  output       io_wt_actv_nz_0_95,
  output       io_wt_actv_nz_0_96,
  output       io_wt_actv_nz_0_97,
  output       io_wt_actv_nz_0_98,
  output       io_wt_actv_nz_0_99,
  output       io_wt_actv_nz_0_100,
  output       io_wt_actv_nz_0_101,
  output       io_wt_actv_nz_0_102,
  output       io_wt_actv_nz_0_103,
  output       io_wt_actv_nz_0_104,
  output       io_wt_actv_nz_0_105,
  output       io_wt_actv_nz_0_106,
  output       io_wt_actv_nz_0_107,
  output       io_wt_actv_nz_0_108,
  output       io_wt_actv_nz_0_109,
  output       io_wt_actv_nz_0_110,
  output       io_wt_actv_nz_0_111,
  output       io_wt_actv_nz_0_112,
  output       io_wt_actv_nz_0_113,
  output       io_wt_actv_nz_0_114,
  output       io_wt_actv_nz_0_115,
  output       io_wt_actv_nz_0_116,
  output       io_wt_actv_nz_0_117,
  output       io_wt_actv_nz_0_118,
  output       io_wt_actv_nz_0_119,
  output       io_wt_actv_nz_0_120,
  output       io_wt_actv_nz_0_121,
  output       io_wt_actv_nz_0_122,
  output       io_wt_actv_nz_0_123,
  output       io_wt_actv_nz_0_124,
  output       io_wt_actv_nz_0_125,
  output       io_wt_actv_nz_0_126,
  output       io_wt_actv_nz_0_127,
  output       io_wt_actv_pvld_0_0,
  output       io_wt_actv_pvld_0_1,
  output       io_wt_actv_pvld_0_2,
  output       io_wt_actv_pvld_0_3,
  output       io_wt_actv_pvld_0_4,
  output       io_wt_actv_pvld_0_5,
  output       io_wt_actv_pvld_0_6,
  output       io_wt_actv_pvld_0_7,
  output       io_wt_actv_pvld_0_8,
  output       io_wt_actv_pvld_0_9,
  output       io_wt_actv_pvld_0_10,
  output       io_wt_actv_pvld_0_11,
  output       io_wt_actv_pvld_0_12,
  output       io_wt_actv_pvld_0_13,
  output       io_wt_actv_pvld_0_14,
  output       io_wt_actv_pvld_0_15,
  output       io_wt_actv_pvld_0_16,
  output       io_wt_actv_pvld_0_17,
  output       io_wt_actv_pvld_0_18,
  output       io_wt_actv_pvld_0_19,
  output       io_wt_actv_pvld_0_20,
  output       io_wt_actv_pvld_0_21,
  output       io_wt_actv_pvld_0_22,
  output       io_wt_actv_pvld_0_23,
  output       io_wt_actv_pvld_0_24,
  output       io_wt_actv_pvld_0_25,
  output       io_wt_actv_pvld_0_26,
  output       io_wt_actv_pvld_0_27,
  output       io_wt_actv_pvld_0_28,
  output       io_wt_actv_pvld_0_29,
  output       io_wt_actv_pvld_0_30,
  output       io_wt_actv_pvld_0_31,
  output       io_wt_actv_pvld_0_32,
  output       io_wt_actv_pvld_0_33,
  output       io_wt_actv_pvld_0_34,
  output       io_wt_actv_pvld_0_35,
  output       io_wt_actv_pvld_0_36,
  output       io_wt_actv_pvld_0_37,
  output       io_wt_actv_pvld_0_38,
  output       io_wt_actv_pvld_0_39,
  output       io_wt_actv_pvld_0_40,
  output       io_wt_actv_pvld_0_41,
  output       io_wt_actv_pvld_0_42,
  output       io_wt_actv_pvld_0_43,
  output       io_wt_actv_pvld_0_44,
  output       io_wt_actv_pvld_0_45,
  output       io_wt_actv_pvld_0_46,
  output       io_wt_actv_pvld_0_47,
  output       io_wt_actv_pvld_0_48,
  output       io_wt_actv_pvld_0_49,
  output       io_wt_actv_pvld_0_50,
  output       io_wt_actv_pvld_0_51,
  output       io_wt_actv_pvld_0_52,
  output       io_wt_actv_pvld_0_53,
  output       io_wt_actv_pvld_0_54,
  output       io_wt_actv_pvld_0_55,
  output       io_wt_actv_pvld_0_56,
  output       io_wt_actv_pvld_0_57,
  output       io_wt_actv_pvld_0_58,
  output       io_wt_actv_pvld_0_59,
  output       io_wt_actv_pvld_0_60,
  output       io_wt_actv_pvld_0_61,
  output       io_wt_actv_pvld_0_62,
  output       io_wt_actv_pvld_0_63,
  output       io_wt_actv_pvld_0_64,
  output       io_wt_actv_pvld_0_65,
  output       io_wt_actv_pvld_0_66,
  output       io_wt_actv_pvld_0_67,
  output       io_wt_actv_pvld_0_68,
  output       io_wt_actv_pvld_0_69,
  output       io_wt_actv_pvld_0_70,
  output       io_wt_actv_pvld_0_71,
  output       io_wt_actv_pvld_0_72,
  output       io_wt_actv_pvld_0_73,
  output       io_wt_actv_pvld_0_74,
  output       io_wt_actv_pvld_0_75,
  output       io_wt_actv_pvld_0_76,
  output       io_wt_actv_pvld_0_77,
  output       io_wt_actv_pvld_0_78,
  output       io_wt_actv_pvld_0_79,
  output       io_wt_actv_pvld_0_80,
  output       io_wt_actv_pvld_0_81,
  output       io_wt_actv_pvld_0_82,
  output       io_wt_actv_pvld_0_83,
  output       io_wt_actv_pvld_0_84,
  output       io_wt_actv_pvld_0_85,
  output       io_wt_actv_pvld_0_86,
  output       io_wt_actv_pvld_0_87,
  output       io_wt_actv_pvld_0_88,
  output       io_wt_actv_pvld_0_89,
  output       io_wt_actv_pvld_0_90,
  output       io_wt_actv_pvld_0_91,
  output       io_wt_actv_pvld_0_92,
  output       io_wt_actv_pvld_0_93,
  output       io_wt_actv_pvld_0_94,
  output       io_wt_actv_pvld_0_95,
  output       io_wt_actv_pvld_0_96,
  output       io_wt_actv_pvld_0_97,
  output       io_wt_actv_pvld_0_98,
  output       io_wt_actv_pvld_0_99,
  output       io_wt_actv_pvld_0_100,
  output       io_wt_actv_pvld_0_101,
  output       io_wt_actv_pvld_0_102,
  output       io_wt_actv_pvld_0_103,
  output       io_wt_actv_pvld_0_104,
  output       io_wt_actv_pvld_0_105,
  output       io_wt_actv_pvld_0_106,
  output       io_wt_actv_pvld_0_107,
  output       io_wt_actv_pvld_0_108,
  output       io_wt_actv_pvld_0_109,
  output       io_wt_actv_pvld_0_110,
  output       io_wt_actv_pvld_0_111,
  output       io_wt_actv_pvld_0_112,
  output       io_wt_actv_pvld_0_113,
  output       io_wt_actv_pvld_0_114,
  output       io_wt_actv_pvld_0_115,
  output       io_wt_actv_pvld_0_116,
  output       io_wt_actv_pvld_0_117,
  output       io_wt_actv_pvld_0_118,
  output       io_wt_actv_pvld_0_119,
  output       io_wt_actv_pvld_0_120,
  output       io_wt_actv_pvld_0_121,
  output       io_wt_actv_pvld_0_122,
  output       io_wt_actv_pvld_0_123,
  output       io_wt_actv_pvld_0_124,
  output       io_wt_actv_pvld_0_125,
  output       io_wt_actv_pvld_0_126,
  output       io_wt_actv_pvld_0_127
);
  reg  wt_pre_nz_0; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_0;
  reg  wt_pre_nz_1; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_1;
  reg  wt_pre_nz_2; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_2;
  reg  wt_pre_nz_3; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_3;
  reg  wt_pre_nz_4; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_4;
  reg  wt_pre_nz_5; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_5;
  reg  wt_pre_nz_6; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_6;
  reg  wt_pre_nz_7; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_7;
  reg  wt_pre_nz_8; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_8;
  reg  wt_pre_nz_9; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_9;
  reg  wt_pre_nz_10; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_10;
  reg  wt_pre_nz_11; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_11;
  reg  wt_pre_nz_12; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_12;
  reg  wt_pre_nz_13; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_13;
  reg  wt_pre_nz_14; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_14;
  reg  wt_pre_nz_15; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_15;
  reg  wt_pre_nz_16; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_16;
  reg  wt_pre_nz_17; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_17;
  reg  wt_pre_nz_18; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_18;
  reg  wt_pre_nz_19; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_19;
  reg  wt_pre_nz_20; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_20;
  reg  wt_pre_nz_21; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_21;
  reg  wt_pre_nz_22; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_22;
  reg  wt_pre_nz_23; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_23;
  reg  wt_pre_nz_24; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_24;
  reg  wt_pre_nz_25; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_25;
  reg  wt_pre_nz_26; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_26;
  reg  wt_pre_nz_27; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_27;
  reg  wt_pre_nz_28; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_28;
  reg  wt_pre_nz_29; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_29;
  reg  wt_pre_nz_30; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_30;
  reg  wt_pre_nz_31; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_31;
  reg  wt_pre_nz_32; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_32;
  reg  wt_pre_nz_33; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_33;
  reg  wt_pre_nz_34; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_34;
  reg  wt_pre_nz_35; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_35;
  reg  wt_pre_nz_36; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_36;
  reg  wt_pre_nz_37; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_37;
  reg  wt_pre_nz_38; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_38;
  reg  wt_pre_nz_39; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_39;
  reg  wt_pre_nz_40; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_40;
  reg  wt_pre_nz_41; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_41;
  reg  wt_pre_nz_42; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_42;
  reg  wt_pre_nz_43; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_43;
  reg  wt_pre_nz_44; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_44;
  reg  wt_pre_nz_45; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_45;
  reg  wt_pre_nz_46; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_46;
  reg  wt_pre_nz_47; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_47;
  reg  wt_pre_nz_48; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_48;
  reg  wt_pre_nz_49; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_49;
  reg  wt_pre_nz_50; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_50;
  reg  wt_pre_nz_51; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_51;
  reg  wt_pre_nz_52; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_52;
  reg  wt_pre_nz_53; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_53;
  reg  wt_pre_nz_54; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_54;
  reg  wt_pre_nz_55; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_55;
  reg  wt_pre_nz_56; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_56;
  reg  wt_pre_nz_57; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_57;
  reg  wt_pre_nz_58; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_58;
  reg  wt_pre_nz_59; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_59;
  reg  wt_pre_nz_60; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_60;
  reg  wt_pre_nz_61; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_61;
  reg  wt_pre_nz_62; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_62;
  reg  wt_pre_nz_63; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_63;
  reg  wt_pre_nz_64; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_64;
  reg  wt_pre_nz_65; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_65;
  reg  wt_pre_nz_66; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_66;
  reg  wt_pre_nz_67; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_67;
  reg  wt_pre_nz_68; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_68;
  reg  wt_pre_nz_69; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_69;
  reg  wt_pre_nz_70; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_70;
  reg  wt_pre_nz_71; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_71;
  reg  wt_pre_nz_72; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_72;
  reg  wt_pre_nz_73; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_73;
  reg  wt_pre_nz_74; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_74;
  reg  wt_pre_nz_75; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_75;
  reg  wt_pre_nz_76; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_76;
  reg  wt_pre_nz_77; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_77;
  reg  wt_pre_nz_78; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_78;
  reg  wt_pre_nz_79; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_79;
  reg  wt_pre_nz_80; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_80;
  reg  wt_pre_nz_81; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_81;
  reg  wt_pre_nz_82; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_82;
  reg  wt_pre_nz_83; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_83;
  reg  wt_pre_nz_84; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_84;
  reg  wt_pre_nz_85; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_85;
  reg  wt_pre_nz_86; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_86;
  reg  wt_pre_nz_87; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_87;
  reg  wt_pre_nz_88; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_88;
  reg  wt_pre_nz_89; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_89;
  reg  wt_pre_nz_90; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_90;
  reg  wt_pre_nz_91; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_91;
  reg  wt_pre_nz_92; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_92;
  reg  wt_pre_nz_93; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_93;
  reg  wt_pre_nz_94; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_94;
  reg  wt_pre_nz_95; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_95;
  reg  wt_pre_nz_96; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_96;
  reg  wt_pre_nz_97; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_97;
  reg  wt_pre_nz_98; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_98;
  reg  wt_pre_nz_99; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_99;
  reg  wt_pre_nz_100; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_100;
  reg  wt_pre_nz_101; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_101;
  reg  wt_pre_nz_102; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_102;
  reg  wt_pre_nz_103; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_103;
  reg  wt_pre_nz_104; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_104;
  reg  wt_pre_nz_105; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_105;
  reg  wt_pre_nz_106; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_106;
  reg  wt_pre_nz_107; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_107;
  reg  wt_pre_nz_108; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_108;
  reg  wt_pre_nz_109; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_109;
  reg  wt_pre_nz_110; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_110;
  reg  wt_pre_nz_111; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_111;
  reg  wt_pre_nz_112; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_112;
  reg  wt_pre_nz_113; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_113;
  reg  wt_pre_nz_114; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_114;
  reg  wt_pre_nz_115; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_115;
  reg  wt_pre_nz_116; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_116;
  reg  wt_pre_nz_117; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_117;
  reg  wt_pre_nz_118; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_118;
  reg  wt_pre_nz_119; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_119;
  reg  wt_pre_nz_120; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_120;
  reg  wt_pre_nz_121; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_121;
  reg  wt_pre_nz_122; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_122;
  reg  wt_pre_nz_123; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_123;
  reg  wt_pre_nz_124; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_124;
  reg  wt_pre_nz_125; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_125;
  reg  wt_pre_nz_126; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_126;
  reg  wt_pre_nz_127; // @[NV_NVDLA_CMAC_CORE_active.scala 65:28]
  reg [31:0] _RAND_127;
  reg [7:0] wt_pre_data_0; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_128;
  reg [7:0] wt_pre_data_1; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_129;
  reg [7:0] wt_pre_data_2; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_130;
  reg [7:0] wt_pre_data_3; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_131;
  reg [7:0] wt_pre_data_4; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_132;
  reg [7:0] wt_pre_data_5; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_133;
  reg [7:0] wt_pre_data_6; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_134;
  reg [7:0] wt_pre_data_7; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_135;
  reg [7:0] wt_pre_data_8; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_136;
  reg [7:0] wt_pre_data_9; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_137;
  reg [7:0] wt_pre_data_10; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_138;
  reg [7:0] wt_pre_data_11; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_139;
  reg [7:0] wt_pre_data_12; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_140;
  reg [7:0] wt_pre_data_13; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_141;
  reg [7:0] wt_pre_data_14; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_142;
  reg [7:0] wt_pre_data_15; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_143;
  reg [7:0] wt_pre_data_16; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_144;
  reg [7:0] wt_pre_data_17; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_145;
  reg [7:0] wt_pre_data_18; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_146;
  reg [7:0] wt_pre_data_19; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_147;
  reg [7:0] wt_pre_data_20; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_148;
  reg [7:0] wt_pre_data_21; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_149;
  reg [7:0] wt_pre_data_22; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_150;
  reg [7:0] wt_pre_data_23; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_151;
  reg [7:0] wt_pre_data_24; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_152;
  reg [7:0] wt_pre_data_25; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_153;
  reg [7:0] wt_pre_data_26; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_154;
  reg [7:0] wt_pre_data_27; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_155;
  reg [7:0] wt_pre_data_28; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_156;
  reg [7:0] wt_pre_data_29; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_157;
  reg [7:0] wt_pre_data_30; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_158;
  reg [7:0] wt_pre_data_31; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_159;
  reg [7:0] wt_pre_data_32; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_160;
  reg [7:0] wt_pre_data_33; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_161;
  reg [7:0] wt_pre_data_34; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_162;
  reg [7:0] wt_pre_data_35; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_163;
  reg [7:0] wt_pre_data_36; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_164;
  reg [7:0] wt_pre_data_37; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_165;
  reg [7:0] wt_pre_data_38; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_166;
  reg [7:0] wt_pre_data_39; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_167;
  reg [7:0] wt_pre_data_40; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_168;
  reg [7:0] wt_pre_data_41; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_169;
  reg [7:0] wt_pre_data_42; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_170;
  reg [7:0] wt_pre_data_43; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_171;
  reg [7:0] wt_pre_data_44; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_172;
  reg [7:0] wt_pre_data_45; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_173;
  reg [7:0] wt_pre_data_46; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_174;
  reg [7:0] wt_pre_data_47; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_175;
  reg [7:0] wt_pre_data_48; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_176;
  reg [7:0] wt_pre_data_49; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_177;
  reg [7:0] wt_pre_data_50; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_178;
  reg [7:0] wt_pre_data_51; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_179;
  reg [7:0] wt_pre_data_52; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_180;
  reg [7:0] wt_pre_data_53; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_181;
  reg [7:0] wt_pre_data_54; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_182;
  reg [7:0] wt_pre_data_55; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_183;
  reg [7:0] wt_pre_data_56; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_184;
  reg [7:0] wt_pre_data_57; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_185;
  reg [7:0] wt_pre_data_58; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_186;
  reg [7:0] wt_pre_data_59; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_187;
  reg [7:0] wt_pre_data_60; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_188;
  reg [7:0] wt_pre_data_61; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_189;
  reg [7:0] wt_pre_data_62; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_190;
  reg [7:0] wt_pre_data_63; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_191;
  reg [7:0] wt_pre_data_64; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_192;
  reg [7:0] wt_pre_data_65; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_193;
  reg [7:0] wt_pre_data_66; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_194;
  reg [7:0] wt_pre_data_67; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_195;
  reg [7:0] wt_pre_data_68; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_196;
  reg [7:0] wt_pre_data_69; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_197;
  reg [7:0] wt_pre_data_70; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_198;
  reg [7:0] wt_pre_data_71; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_199;
  reg [7:0] wt_pre_data_72; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_200;
  reg [7:0] wt_pre_data_73; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_201;
  reg [7:0] wt_pre_data_74; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_202;
  reg [7:0] wt_pre_data_75; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_203;
  reg [7:0] wt_pre_data_76; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_204;
  reg [7:0] wt_pre_data_77; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_205;
  reg [7:0] wt_pre_data_78; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_206;
  reg [7:0] wt_pre_data_79; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_207;
  reg [7:0] wt_pre_data_80; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_208;
  reg [7:0] wt_pre_data_81; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_209;
  reg [7:0] wt_pre_data_82; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_210;
  reg [7:0] wt_pre_data_83; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_211;
  reg [7:0] wt_pre_data_84; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_212;
  reg [7:0] wt_pre_data_85; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_213;
  reg [7:0] wt_pre_data_86; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_214;
  reg [7:0] wt_pre_data_87; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_215;
  reg [7:0] wt_pre_data_88; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_216;
  reg [7:0] wt_pre_data_89; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_217;
  reg [7:0] wt_pre_data_90; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_218;
  reg [7:0] wt_pre_data_91; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_219;
  reg [7:0] wt_pre_data_92; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_220;
  reg [7:0] wt_pre_data_93; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_221;
  reg [7:0] wt_pre_data_94; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_222;
  reg [7:0] wt_pre_data_95; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_223;
  reg [7:0] wt_pre_data_96; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_224;
  reg [7:0] wt_pre_data_97; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_225;
  reg [7:0] wt_pre_data_98; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_226;
  reg [7:0] wt_pre_data_99; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_227;
  reg [7:0] wt_pre_data_100; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_228;
  reg [7:0] wt_pre_data_101; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_229;
  reg [7:0] wt_pre_data_102; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_230;
  reg [7:0] wt_pre_data_103; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_231;
  reg [7:0] wt_pre_data_104; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_232;
  reg [7:0] wt_pre_data_105; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_233;
  reg [7:0] wt_pre_data_106; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_234;
  reg [7:0] wt_pre_data_107; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_235;
  reg [7:0] wt_pre_data_108; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_236;
  reg [7:0] wt_pre_data_109; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_237;
  reg [7:0] wt_pre_data_110; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_238;
  reg [7:0] wt_pre_data_111; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_239;
  reg [7:0] wt_pre_data_112; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_240;
  reg [7:0] wt_pre_data_113; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_241;
  reg [7:0] wt_pre_data_114; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_242;
  reg [7:0] wt_pre_data_115; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_243;
  reg [7:0] wt_pre_data_116; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_244;
  reg [7:0] wt_pre_data_117; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_245;
  reg [7:0] wt_pre_data_118; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_246;
  reg [7:0] wt_pre_data_119; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_247;
  reg [7:0] wt_pre_data_120; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_248;
  reg [7:0] wt_pre_data_121; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_249;
  reg [7:0] wt_pre_data_122; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_250;
  reg [7:0] wt_pre_data_123; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_251;
  reg [7:0] wt_pre_data_124; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_252;
  reg [7:0] wt_pre_data_125; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_253;
  reg [7:0] wt_pre_data_126; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_254;
  reg [7:0] wt_pre_data_127; // @[NV_NVDLA_CMAC_CORE_active.scala 66:26]
  reg [31:0] _RAND_255;
  reg  wt_pre_sel_0; // @[NV_NVDLA_CMAC_CORE_active.scala 67:29]
  reg [31:0] _RAND_256;
  wire [7:0] _GEN_0; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_1; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_2; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_3; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_4; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_5; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_6; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_7; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_8; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_9; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_10; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_11; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_12; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_13; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_14; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_15; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_16; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_17; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_18; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_19; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_20; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_21; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_22; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_23; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_24; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_25; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_26; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_27; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_28; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_29; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_30; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_31; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_32; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_33; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_34; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_35; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_36; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_37; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_38; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_39; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_40; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_41; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_42; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_43; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_44; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_45; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_46; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_47; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_48; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_49; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_50; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_51; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_52; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_53; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_54; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_55; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_56; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_57; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_58; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_59; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_60; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_61; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_62; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_63; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_64; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_65; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_66; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_67; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_68; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_69; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_70; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_71; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_72; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_73; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_74; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_75; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_76; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_77; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_78; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_79; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_80; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_81; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_82; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_83; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_84; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_85; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_86; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_87; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_88; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_89; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_90; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_91; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_92; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_93; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_94; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_95; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_96; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_97; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_98; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_99; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_100; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_101; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_102; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_103; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_104; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_105; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_106; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_107; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_108; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_109; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_110; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_111; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_112; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_113; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_114; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_115; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_116; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_117; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_118; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_119; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_120; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_121; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_122; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_123; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_124; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_125; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_126; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire [7:0] _GEN_127; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  wire  _GEN_128; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_129; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_130; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_131; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_132; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_133; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_134; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_135; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_136; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_137; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_138; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_139; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_140; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_141; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_142; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_143; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_144; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_145; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_146; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_147; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_148; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_149; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_150; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_151; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_152; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_153; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_154; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_155; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_156; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_157; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_158; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_159; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_160; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_161; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_162; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_163; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_164; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_165; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_166; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_167; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_168; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_169; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_170; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_171; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_172; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_173; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_174; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_175; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_176; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_177; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_178; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_179; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_180; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_181; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_182; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_183; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_184; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_185; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_186; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_187; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_188; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_189; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_190; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_191; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_192; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_193; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_194; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_195; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_196; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_197; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_198; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_199; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_200; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_201; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_202; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_203; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_204; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_205; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_206; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_207; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_208; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_209; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_210; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_211; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_212; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_213; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_214; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_215; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_216; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_217; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_218; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_219; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_220; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_221; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_222; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_223; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_224; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_225; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_226; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_227; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_228; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_229; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_230; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_231; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_232; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_233; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_234; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_235; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_236; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_237; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_238; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_239; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_240; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_241; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_242; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_243; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_244; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_245; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_246; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_247; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_248; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_249; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_250; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_251; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_252; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_253; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_254; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_255; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  wire  _GEN_256; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  reg  dat_pre_nz_0; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_257;
  reg  dat_pre_nz_1; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_258;
  reg  dat_pre_nz_2; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_259;
  reg  dat_pre_nz_3; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_260;
  reg  dat_pre_nz_4; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_261;
  reg  dat_pre_nz_5; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_262;
  reg  dat_pre_nz_6; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_263;
  reg  dat_pre_nz_7; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_264;
  reg  dat_pre_nz_8; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_265;
  reg  dat_pre_nz_9; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_266;
  reg  dat_pre_nz_10; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_267;
  reg  dat_pre_nz_11; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_268;
  reg  dat_pre_nz_12; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_269;
  reg  dat_pre_nz_13; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_270;
  reg  dat_pre_nz_14; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_271;
  reg  dat_pre_nz_15; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_272;
  reg  dat_pre_nz_16; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_273;
  reg  dat_pre_nz_17; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_274;
  reg  dat_pre_nz_18; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_275;
  reg  dat_pre_nz_19; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_276;
  reg  dat_pre_nz_20; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_277;
  reg  dat_pre_nz_21; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_278;
  reg  dat_pre_nz_22; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_279;
  reg  dat_pre_nz_23; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_280;
  reg  dat_pre_nz_24; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_281;
  reg  dat_pre_nz_25; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_282;
  reg  dat_pre_nz_26; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_283;
  reg  dat_pre_nz_27; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_284;
  reg  dat_pre_nz_28; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_285;
  reg  dat_pre_nz_29; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_286;
  reg  dat_pre_nz_30; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_287;
  reg  dat_pre_nz_31; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_288;
  reg  dat_pre_nz_32; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_289;
  reg  dat_pre_nz_33; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_290;
  reg  dat_pre_nz_34; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_291;
  reg  dat_pre_nz_35; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_292;
  reg  dat_pre_nz_36; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_293;
  reg  dat_pre_nz_37; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_294;
  reg  dat_pre_nz_38; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_295;
  reg  dat_pre_nz_39; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_296;
  reg  dat_pre_nz_40; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_297;
  reg  dat_pre_nz_41; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_298;
  reg  dat_pre_nz_42; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_299;
  reg  dat_pre_nz_43; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_300;
  reg  dat_pre_nz_44; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_301;
  reg  dat_pre_nz_45; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_302;
  reg  dat_pre_nz_46; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_303;
  reg  dat_pre_nz_47; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_304;
  reg  dat_pre_nz_48; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_305;
  reg  dat_pre_nz_49; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_306;
  reg  dat_pre_nz_50; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_307;
  reg  dat_pre_nz_51; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_308;
  reg  dat_pre_nz_52; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_309;
  reg  dat_pre_nz_53; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_310;
  reg  dat_pre_nz_54; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_311;
  reg  dat_pre_nz_55; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_312;
  reg  dat_pre_nz_56; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_313;
  reg  dat_pre_nz_57; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_314;
  reg  dat_pre_nz_58; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_315;
  reg  dat_pre_nz_59; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_316;
  reg  dat_pre_nz_60; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_317;
  reg  dat_pre_nz_61; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_318;
  reg  dat_pre_nz_62; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_319;
  reg  dat_pre_nz_63; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_320;
  reg  dat_pre_nz_64; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_321;
  reg  dat_pre_nz_65; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_322;
  reg  dat_pre_nz_66; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_323;
  reg  dat_pre_nz_67; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_324;
  reg  dat_pre_nz_68; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_325;
  reg  dat_pre_nz_69; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_326;
  reg  dat_pre_nz_70; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_327;
  reg  dat_pre_nz_71; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_328;
  reg  dat_pre_nz_72; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_329;
  reg  dat_pre_nz_73; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_330;
  reg  dat_pre_nz_74; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_331;
  reg  dat_pre_nz_75; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_332;
  reg  dat_pre_nz_76; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_333;
  reg  dat_pre_nz_77; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_334;
  reg  dat_pre_nz_78; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_335;
  reg  dat_pre_nz_79; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_336;
  reg  dat_pre_nz_80; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_337;
  reg  dat_pre_nz_81; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_338;
  reg  dat_pre_nz_82; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_339;
  reg  dat_pre_nz_83; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_340;
  reg  dat_pre_nz_84; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_341;
  reg  dat_pre_nz_85; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_342;
  reg  dat_pre_nz_86; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_343;
  reg  dat_pre_nz_87; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_344;
  reg  dat_pre_nz_88; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_345;
  reg  dat_pre_nz_89; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_346;
  reg  dat_pre_nz_90; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_347;
  reg  dat_pre_nz_91; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_348;
  reg  dat_pre_nz_92; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_349;
  reg  dat_pre_nz_93; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_350;
  reg  dat_pre_nz_94; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_351;
  reg  dat_pre_nz_95; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_352;
  reg  dat_pre_nz_96; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_353;
  reg  dat_pre_nz_97; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_354;
  reg  dat_pre_nz_98; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_355;
  reg  dat_pre_nz_99; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_356;
  reg  dat_pre_nz_100; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_357;
  reg  dat_pre_nz_101; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_358;
  reg  dat_pre_nz_102; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_359;
  reg  dat_pre_nz_103; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_360;
  reg  dat_pre_nz_104; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_361;
  reg  dat_pre_nz_105; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_362;
  reg  dat_pre_nz_106; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_363;
  reg  dat_pre_nz_107; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_364;
  reg  dat_pre_nz_108; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_365;
  reg  dat_pre_nz_109; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_366;
  reg  dat_pre_nz_110; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_367;
  reg  dat_pre_nz_111; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_368;
  reg  dat_pre_nz_112; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_369;
  reg  dat_pre_nz_113; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_370;
  reg  dat_pre_nz_114; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_371;
  reg  dat_pre_nz_115; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_372;
  reg  dat_pre_nz_116; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_373;
  reg  dat_pre_nz_117; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_374;
  reg  dat_pre_nz_118; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_375;
  reg  dat_pre_nz_119; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_376;
  reg  dat_pre_nz_120; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_377;
  reg  dat_pre_nz_121; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_378;
  reg  dat_pre_nz_122; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_379;
  reg  dat_pre_nz_123; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_380;
  reg  dat_pre_nz_124; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_381;
  reg  dat_pre_nz_125; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_382;
  reg  dat_pre_nz_126; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_383;
  reg  dat_pre_nz_127; // @[NV_NVDLA_CMAC_CORE_active.scala 82:29]
  reg [31:0] _RAND_384;
  reg [7:0] dat_pre_data_0; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_385;
  reg [7:0] dat_pre_data_1; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_386;
  reg [7:0] dat_pre_data_2; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_387;
  reg [7:0] dat_pre_data_3; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_388;
  reg [7:0] dat_pre_data_4; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_389;
  reg [7:0] dat_pre_data_5; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_390;
  reg [7:0] dat_pre_data_6; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_391;
  reg [7:0] dat_pre_data_7; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_392;
  reg [7:0] dat_pre_data_8; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_393;
  reg [7:0] dat_pre_data_9; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_394;
  reg [7:0] dat_pre_data_10; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_395;
  reg [7:0] dat_pre_data_11; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_396;
  reg [7:0] dat_pre_data_12; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_397;
  reg [7:0] dat_pre_data_13; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_398;
  reg [7:0] dat_pre_data_14; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_399;
  reg [7:0] dat_pre_data_15; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_400;
  reg [7:0] dat_pre_data_16; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_401;
  reg [7:0] dat_pre_data_17; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_402;
  reg [7:0] dat_pre_data_18; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_403;
  reg [7:0] dat_pre_data_19; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_404;
  reg [7:0] dat_pre_data_20; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_405;
  reg [7:0] dat_pre_data_21; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_406;
  reg [7:0] dat_pre_data_22; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_407;
  reg [7:0] dat_pre_data_23; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_408;
  reg [7:0] dat_pre_data_24; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_409;
  reg [7:0] dat_pre_data_25; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_410;
  reg [7:0] dat_pre_data_26; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_411;
  reg [7:0] dat_pre_data_27; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_412;
  reg [7:0] dat_pre_data_28; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_413;
  reg [7:0] dat_pre_data_29; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_414;
  reg [7:0] dat_pre_data_30; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_415;
  reg [7:0] dat_pre_data_31; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_416;
  reg [7:0] dat_pre_data_32; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_417;
  reg [7:0] dat_pre_data_33; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_418;
  reg [7:0] dat_pre_data_34; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_419;
  reg [7:0] dat_pre_data_35; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_420;
  reg [7:0] dat_pre_data_36; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_421;
  reg [7:0] dat_pre_data_37; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_422;
  reg [7:0] dat_pre_data_38; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_423;
  reg [7:0] dat_pre_data_39; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_424;
  reg [7:0] dat_pre_data_40; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_425;
  reg [7:0] dat_pre_data_41; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_426;
  reg [7:0] dat_pre_data_42; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_427;
  reg [7:0] dat_pre_data_43; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_428;
  reg [7:0] dat_pre_data_44; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_429;
  reg [7:0] dat_pre_data_45; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_430;
  reg [7:0] dat_pre_data_46; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_431;
  reg [7:0] dat_pre_data_47; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_432;
  reg [7:0] dat_pre_data_48; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_433;
  reg [7:0] dat_pre_data_49; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_434;
  reg [7:0] dat_pre_data_50; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_435;
  reg [7:0] dat_pre_data_51; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_436;
  reg [7:0] dat_pre_data_52; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_437;
  reg [7:0] dat_pre_data_53; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_438;
  reg [7:0] dat_pre_data_54; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_439;
  reg [7:0] dat_pre_data_55; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_440;
  reg [7:0] dat_pre_data_56; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_441;
  reg [7:0] dat_pre_data_57; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_442;
  reg [7:0] dat_pre_data_58; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_443;
  reg [7:0] dat_pre_data_59; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_444;
  reg [7:0] dat_pre_data_60; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_445;
  reg [7:0] dat_pre_data_61; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_446;
  reg [7:0] dat_pre_data_62; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_447;
  reg [7:0] dat_pre_data_63; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_448;
  reg [7:0] dat_pre_data_64; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_449;
  reg [7:0] dat_pre_data_65; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_450;
  reg [7:0] dat_pre_data_66; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_451;
  reg [7:0] dat_pre_data_67; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_452;
  reg [7:0] dat_pre_data_68; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_453;
  reg [7:0] dat_pre_data_69; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_454;
  reg [7:0] dat_pre_data_70; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_455;
  reg [7:0] dat_pre_data_71; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_456;
  reg [7:0] dat_pre_data_72; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_457;
  reg [7:0] dat_pre_data_73; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_458;
  reg [7:0] dat_pre_data_74; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_459;
  reg [7:0] dat_pre_data_75; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_460;
  reg [7:0] dat_pre_data_76; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_461;
  reg [7:0] dat_pre_data_77; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_462;
  reg [7:0] dat_pre_data_78; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_463;
  reg [7:0] dat_pre_data_79; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_464;
  reg [7:0] dat_pre_data_80; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_465;
  reg [7:0] dat_pre_data_81; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_466;
  reg [7:0] dat_pre_data_82; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_467;
  reg [7:0] dat_pre_data_83; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_468;
  reg [7:0] dat_pre_data_84; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_469;
  reg [7:0] dat_pre_data_85; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_470;
  reg [7:0] dat_pre_data_86; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_471;
  reg [7:0] dat_pre_data_87; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_472;
  reg [7:0] dat_pre_data_88; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_473;
  reg [7:0] dat_pre_data_89; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_474;
  reg [7:0] dat_pre_data_90; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_475;
  reg [7:0] dat_pre_data_91; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_476;
  reg [7:0] dat_pre_data_92; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_477;
  reg [7:0] dat_pre_data_93; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_478;
  reg [7:0] dat_pre_data_94; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_479;
  reg [7:0] dat_pre_data_95; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_480;
  reg [7:0] dat_pre_data_96; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_481;
  reg [7:0] dat_pre_data_97; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_482;
  reg [7:0] dat_pre_data_98; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_483;
  reg [7:0] dat_pre_data_99; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_484;
  reg [7:0] dat_pre_data_100; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_485;
  reg [7:0] dat_pre_data_101; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_486;
  reg [7:0] dat_pre_data_102; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_487;
  reg [7:0] dat_pre_data_103; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_488;
  reg [7:0] dat_pre_data_104; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_489;
  reg [7:0] dat_pre_data_105; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_490;
  reg [7:0] dat_pre_data_106; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_491;
  reg [7:0] dat_pre_data_107; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_492;
  reg [7:0] dat_pre_data_108; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_493;
  reg [7:0] dat_pre_data_109; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_494;
  reg [7:0] dat_pre_data_110; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_495;
  reg [7:0] dat_pre_data_111; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_496;
  reg [7:0] dat_pre_data_112; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_497;
  reg [7:0] dat_pre_data_113; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_498;
  reg [7:0] dat_pre_data_114; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_499;
  reg [7:0] dat_pre_data_115; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_500;
  reg [7:0] dat_pre_data_116; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_501;
  reg [7:0] dat_pre_data_117; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_502;
  reg [7:0] dat_pre_data_118; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_503;
  reg [7:0] dat_pre_data_119; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_504;
  reg [7:0] dat_pre_data_120; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_505;
  reg [7:0] dat_pre_data_121; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_506;
  reg [7:0] dat_pre_data_122; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_507;
  reg [7:0] dat_pre_data_123; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_508;
  reg [7:0] dat_pre_data_124; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_509;
  reg [7:0] dat_pre_data_125; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_510;
  reg [7:0] dat_pre_data_126; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_511;
  reg [7:0] dat_pre_data_127; // @[NV_NVDLA_CMAC_CORE_active.scala 83:27]
  reg [31:0] _RAND_512;
  reg  dat_pre_pvld; // @[NV_NVDLA_CMAC_CORE_active.scala 84:31]
  reg [31:0] _RAND_513;
  reg  dat_pre_stripe_st_out_0; // @[NV_NVDLA_CMAC_CORE_active.scala 85:40]
  reg [31:0] _RAND_514;
  reg  dat_pre_stripe_end_out_0; // @[NV_NVDLA_CMAC_CORE_active.scala 86:41]
  reg [31:0] _RAND_515;
  wire [7:0] _GEN_385; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_386; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_387; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_388; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_389; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_390; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_391; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_392; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_393; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_394; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_395; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_396; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_397; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_398; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_399; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_400; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_401; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_402; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_403; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_404; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_405; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_406; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_407; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_408; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_409; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_410; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_411; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_412; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_413; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_414; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_415; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_416; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_417; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_418; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_419; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_420; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_421; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_422; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_423; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_424; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_425; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_426; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_427; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_428; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_429; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_430; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_431; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_432; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_433; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_434; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_435; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_436; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_437; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_438; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_439; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_440; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_441; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_442; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_443; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_444; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_445; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_446; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_447; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_448; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_449; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_450; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_451; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_452; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_453; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_454; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_455; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_456; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_457; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_458; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_459; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_460; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_461; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_462; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_463; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_464; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_465; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_466; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_467; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_468; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_469; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_470; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_471; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_472; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_473; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_474; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_475; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_476; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_477; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_478; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_479; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_480; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_481; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_482; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_483; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_484; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_485; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_486; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_487; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_488; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_489; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_490; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_491; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_492; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_493; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_494; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_495; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_496; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_497; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_498; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_499; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_500; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_501; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_502; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_503; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_504; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_505; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_506; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_507; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_508; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_509; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_510; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_511; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire [7:0] _GEN_512; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  wire  _GEN_513; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_514; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_515; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_516; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_517; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_518; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_519; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_520; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_521; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_522; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_523; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_524; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_525; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_526; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_527; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_528; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_529; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_530; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_531; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_532; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_533; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_534; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_535; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_536; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_537; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_538; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_539; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_540; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_541; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_542; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_543; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_544; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_545; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_546; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_547; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_548; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_549; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_550; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_551; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_552; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_553; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_554; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_555; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_556; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_557; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_558; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_559; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_560; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_561; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_562; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_563; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_564; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_565; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_566; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_567; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_568; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_569; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_570; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_571; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_572; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_573; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_574; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_575; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_576; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_577; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_578; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_579; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_580; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_581; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_582; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_583; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_584; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_585; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_586; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_587; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_588; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_589; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_590; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_591; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_592; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_593; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_594; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_595; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_596; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_597; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_598; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_599; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_600; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_601; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_602; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_603; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_604; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_605; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_606; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_607; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_608; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_609; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_610; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_611; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_612; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_613; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_614; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_615; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_616; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_617; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_618; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_619; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_620; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_621; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_622; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_623; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_624; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_625; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_626; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_627; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_628; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_629; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_630; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_631; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_632; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_633; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_634; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_635; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_636; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_637; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_638; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_639; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_640; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_769; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  wire  _GEN_770; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  reg  wt_sd_pvld_0; // @[NV_NVDLA_CMAC_CORE_active.scala 108:29]
  reg [31:0] _RAND_516;
  reg  wt_sd_nz_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_517;
  reg  wt_sd_nz_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_518;
  reg  wt_sd_nz_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_519;
  reg  wt_sd_nz_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_520;
  reg  wt_sd_nz_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_521;
  reg  wt_sd_nz_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_522;
  reg  wt_sd_nz_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_523;
  reg  wt_sd_nz_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_524;
  reg  wt_sd_nz_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_525;
  reg  wt_sd_nz_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_526;
  reg  wt_sd_nz_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_527;
  reg  wt_sd_nz_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_528;
  reg  wt_sd_nz_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_529;
  reg  wt_sd_nz_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_530;
  reg  wt_sd_nz_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_531;
  reg  wt_sd_nz_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_532;
  reg  wt_sd_nz_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_533;
  reg  wt_sd_nz_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_534;
  reg  wt_sd_nz_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_535;
  reg  wt_sd_nz_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_536;
  reg  wt_sd_nz_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_537;
  reg  wt_sd_nz_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_538;
  reg  wt_sd_nz_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_539;
  reg  wt_sd_nz_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_540;
  reg  wt_sd_nz_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_541;
  reg  wt_sd_nz_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_542;
  reg  wt_sd_nz_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_543;
  reg  wt_sd_nz_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_544;
  reg  wt_sd_nz_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_545;
  reg  wt_sd_nz_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_546;
  reg  wt_sd_nz_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_547;
  reg  wt_sd_nz_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_548;
  reg  wt_sd_nz_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_549;
  reg  wt_sd_nz_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_550;
  reg  wt_sd_nz_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_551;
  reg  wt_sd_nz_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_552;
  reg  wt_sd_nz_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_553;
  reg  wt_sd_nz_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_554;
  reg  wt_sd_nz_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_555;
  reg  wt_sd_nz_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_556;
  reg  wt_sd_nz_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_557;
  reg  wt_sd_nz_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_558;
  reg  wt_sd_nz_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_559;
  reg  wt_sd_nz_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_560;
  reg  wt_sd_nz_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_561;
  reg  wt_sd_nz_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_562;
  reg  wt_sd_nz_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_563;
  reg  wt_sd_nz_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_564;
  reg  wt_sd_nz_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_565;
  reg  wt_sd_nz_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_566;
  reg  wt_sd_nz_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_567;
  reg  wt_sd_nz_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_568;
  reg  wt_sd_nz_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_569;
  reg  wt_sd_nz_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_570;
  reg  wt_sd_nz_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_571;
  reg  wt_sd_nz_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_572;
  reg  wt_sd_nz_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_573;
  reg  wt_sd_nz_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_574;
  reg  wt_sd_nz_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_575;
  reg  wt_sd_nz_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_576;
  reg  wt_sd_nz_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_577;
  reg  wt_sd_nz_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_578;
  reg  wt_sd_nz_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_579;
  reg  wt_sd_nz_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_580;
  reg  wt_sd_nz_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_581;
  reg  wt_sd_nz_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_582;
  reg  wt_sd_nz_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_583;
  reg  wt_sd_nz_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_584;
  reg  wt_sd_nz_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_585;
  reg  wt_sd_nz_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_586;
  reg  wt_sd_nz_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_587;
  reg  wt_sd_nz_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_588;
  reg  wt_sd_nz_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_589;
  reg  wt_sd_nz_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_590;
  reg  wt_sd_nz_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_591;
  reg  wt_sd_nz_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_592;
  reg  wt_sd_nz_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_593;
  reg  wt_sd_nz_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_594;
  reg  wt_sd_nz_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_595;
  reg  wt_sd_nz_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_596;
  reg  wt_sd_nz_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_597;
  reg  wt_sd_nz_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_598;
  reg  wt_sd_nz_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_599;
  reg  wt_sd_nz_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_600;
  reg  wt_sd_nz_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_601;
  reg  wt_sd_nz_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_602;
  reg  wt_sd_nz_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_603;
  reg  wt_sd_nz_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_604;
  reg  wt_sd_nz_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_605;
  reg  wt_sd_nz_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_606;
  reg  wt_sd_nz_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_607;
  reg  wt_sd_nz_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_608;
  reg  wt_sd_nz_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_609;
  reg  wt_sd_nz_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_610;
  reg  wt_sd_nz_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_611;
  reg  wt_sd_nz_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_612;
  reg  wt_sd_nz_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_613;
  reg  wt_sd_nz_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_614;
  reg  wt_sd_nz_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_615;
  reg  wt_sd_nz_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_616;
  reg  wt_sd_nz_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_617;
  reg  wt_sd_nz_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_618;
  reg  wt_sd_nz_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_619;
  reg  wt_sd_nz_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_620;
  reg  wt_sd_nz_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_621;
  reg  wt_sd_nz_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_622;
  reg  wt_sd_nz_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_623;
  reg  wt_sd_nz_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_624;
  reg  wt_sd_nz_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_625;
  reg  wt_sd_nz_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_626;
  reg  wt_sd_nz_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_627;
  reg  wt_sd_nz_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_628;
  reg  wt_sd_nz_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_629;
  reg  wt_sd_nz_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_630;
  reg  wt_sd_nz_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_631;
  reg  wt_sd_nz_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_632;
  reg  wt_sd_nz_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_633;
  reg  wt_sd_nz_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_634;
  reg  wt_sd_nz_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_635;
  reg  wt_sd_nz_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_636;
  reg  wt_sd_nz_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_637;
  reg  wt_sd_nz_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_638;
  reg  wt_sd_nz_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_639;
  reg  wt_sd_nz_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_640;
  reg  wt_sd_nz_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_641;
  reg  wt_sd_nz_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_642;
  reg  wt_sd_nz_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_643;
  reg  wt_sd_nz_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 110:27]
  reg [31:0] _RAND_644;
  reg [7:0] wt_sd_data_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_645;
  reg [7:0] wt_sd_data_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_646;
  reg [7:0] wt_sd_data_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_647;
  reg [7:0] wt_sd_data_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_648;
  reg [7:0] wt_sd_data_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_649;
  reg [7:0] wt_sd_data_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_650;
  reg [7:0] wt_sd_data_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_651;
  reg [7:0] wt_sd_data_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_652;
  reg [7:0] wt_sd_data_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_653;
  reg [7:0] wt_sd_data_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_654;
  reg [7:0] wt_sd_data_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_655;
  reg [7:0] wt_sd_data_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_656;
  reg [7:0] wt_sd_data_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_657;
  reg [7:0] wt_sd_data_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_658;
  reg [7:0] wt_sd_data_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_659;
  reg [7:0] wt_sd_data_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_660;
  reg [7:0] wt_sd_data_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_661;
  reg [7:0] wt_sd_data_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_662;
  reg [7:0] wt_sd_data_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_663;
  reg [7:0] wt_sd_data_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_664;
  reg [7:0] wt_sd_data_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_665;
  reg [7:0] wt_sd_data_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_666;
  reg [7:0] wt_sd_data_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_667;
  reg [7:0] wt_sd_data_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_668;
  reg [7:0] wt_sd_data_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_669;
  reg [7:0] wt_sd_data_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_670;
  reg [7:0] wt_sd_data_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_671;
  reg [7:0] wt_sd_data_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_672;
  reg [7:0] wt_sd_data_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_673;
  reg [7:0] wt_sd_data_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_674;
  reg [7:0] wt_sd_data_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_675;
  reg [7:0] wt_sd_data_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_676;
  reg [7:0] wt_sd_data_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_677;
  reg [7:0] wt_sd_data_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_678;
  reg [7:0] wt_sd_data_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_679;
  reg [7:0] wt_sd_data_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_680;
  reg [7:0] wt_sd_data_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_681;
  reg [7:0] wt_sd_data_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_682;
  reg [7:0] wt_sd_data_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_683;
  reg [7:0] wt_sd_data_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_684;
  reg [7:0] wt_sd_data_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_685;
  reg [7:0] wt_sd_data_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_686;
  reg [7:0] wt_sd_data_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_687;
  reg [7:0] wt_sd_data_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_688;
  reg [7:0] wt_sd_data_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_689;
  reg [7:0] wt_sd_data_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_690;
  reg [7:0] wt_sd_data_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_691;
  reg [7:0] wt_sd_data_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_692;
  reg [7:0] wt_sd_data_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_693;
  reg [7:0] wt_sd_data_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_694;
  reg [7:0] wt_sd_data_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_695;
  reg [7:0] wt_sd_data_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_696;
  reg [7:0] wt_sd_data_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_697;
  reg [7:0] wt_sd_data_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_698;
  reg [7:0] wt_sd_data_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_699;
  reg [7:0] wt_sd_data_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_700;
  reg [7:0] wt_sd_data_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_701;
  reg [7:0] wt_sd_data_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_702;
  reg [7:0] wt_sd_data_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_703;
  reg [7:0] wt_sd_data_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_704;
  reg [7:0] wt_sd_data_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_705;
  reg [7:0] wt_sd_data_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_706;
  reg [7:0] wt_sd_data_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_707;
  reg [7:0] wt_sd_data_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_708;
  reg [7:0] wt_sd_data_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_709;
  reg [7:0] wt_sd_data_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_710;
  reg [7:0] wt_sd_data_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_711;
  reg [7:0] wt_sd_data_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_712;
  reg [7:0] wt_sd_data_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_713;
  reg [7:0] wt_sd_data_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_714;
  reg [7:0] wt_sd_data_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_715;
  reg [7:0] wt_sd_data_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_716;
  reg [7:0] wt_sd_data_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_717;
  reg [7:0] wt_sd_data_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_718;
  reg [7:0] wt_sd_data_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_719;
  reg [7:0] wt_sd_data_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_720;
  reg [7:0] wt_sd_data_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_721;
  reg [7:0] wt_sd_data_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_722;
  reg [7:0] wt_sd_data_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_723;
  reg [7:0] wt_sd_data_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_724;
  reg [7:0] wt_sd_data_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_725;
  reg [7:0] wt_sd_data_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_726;
  reg [7:0] wt_sd_data_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_727;
  reg [7:0] wt_sd_data_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_728;
  reg [7:0] wt_sd_data_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_729;
  reg [7:0] wt_sd_data_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_730;
  reg [7:0] wt_sd_data_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_731;
  reg [7:0] wt_sd_data_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_732;
  reg [7:0] wt_sd_data_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_733;
  reg [7:0] wt_sd_data_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_734;
  reg [7:0] wt_sd_data_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_735;
  reg [7:0] wt_sd_data_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_736;
  reg [7:0] wt_sd_data_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_737;
  reg [7:0] wt_sd_data_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_738;
  reg [7:0] wt_sd_data_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_739;
  reg [7:0] wt_sd_data_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_740;
  reg [7:0] wt_sd_data_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_741;
  reg [7:0] wt_sd_data_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_742;
  reg [7:0] wt_sd_data_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_743;
  reg [7:0] wt_sd_data_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_744;
  reg [7:0] wt_sd_data_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_745;
  reg [7:0] wt_sd_data_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_746;
  reg [7:0] wt_sd_data_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_747;
  reg [7:0] wt_sd_data_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_748;
  reg [7:0] wt_sd_data_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_749;
  reg [7:0] wt_sd_data_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_750;
  reg [7:0] wt_sd_data_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_751;
  reg [7:0] wt_sd_data_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_752;
  reg [7:0] wt_sd_data_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_753;
  reg [7:0] wt_sd_data_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_754;
  reg [7:0] wt_sd_data_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_755;
  reg [7:0] wt_sd_data_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_756;
  reg [7:0] wt_sd_data_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_757;
  reg [7:0] wt_sd_data_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_758;
  reg [7:0] wt_sd_data_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_759;
  reg [7:0] wt_sd_data_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_760;
  reg [7:0] wt_sd_data_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_761;
  reg [7:0] wt_sd_data_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_762;
  reg [7:0] wt_sd_data_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_763;
  reg [7:0] wt_sd_data_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_764;
  reg [7:0] wt_sd_data_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_765;
  reg [7:0] wt_sd_data_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_766;
  reg [7:0] wt_sd_data_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_767;
  reg [7:0] wt_sd_data_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_768;
  reg [7:0] wt_sd_data_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_769;
  reg [7:0] wt_sd_data_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_770;
  reg [7:0] wt_sd_data_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_771;
  reg [7:0] wt_sd_data_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 111:25]
  reg [31:0] _RAND_772;
  reg  dat_actv_stripe_end_0; // @[NV_NVDLA_CMAC_CORE_active.scala 112:38]
  reg [31:0] _RAND_773;
  wire  _T_27793; // @[NV_NVDLA_CMAC_CORE_active.scala 115:58]
  wire  wt_sd_pvld_w_0; // @[NV_NVDLA_CMAC_CORE_active.scala 115:31]
  wire [7:0] _GEN_771; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_772; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_773; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_774; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_775; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_776; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_777; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_778; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_779; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_780; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_781; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_782; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_783; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_784; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_785; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_786; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_787; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_788; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_789; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_790; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_791; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_792; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_793; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_794; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_795; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_796; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_797; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_798; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_799; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_800; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_801; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_802; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_803; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_804; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_805; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_806; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_807; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_808; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_809; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_810; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_811; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_812; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_813; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_814; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_815; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_816; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_817; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_818; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_819; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_820; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_821; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_822; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_823; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_824; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_825; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_826; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_827; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_828; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_829; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_830; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_831; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_832; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_833; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_834; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_835; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_836; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_837; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_838; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_839; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_840; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_841; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_842; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_843; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_844; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_845; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_846; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_847; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_848; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_849; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_850; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_851; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_852; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_853; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_854; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_855; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_856; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_857; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_858; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_859; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_860; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_861; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_862; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_863; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_864; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_865; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_866; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_867; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_868; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_869; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_870; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_871; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_872; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_873; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_874; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_875; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_876; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_877; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_878; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_879; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_880; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_881; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_882; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_883; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_884; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_885; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_886; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_887; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_888; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_889; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_890; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_891; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_892; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_893; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_894; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_895; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_896; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_897; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire [7:0] _GEN_898; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  wire  _GEN_899; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_900; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_901; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_902; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_903; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_904; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_905; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_906; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_907; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_908; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_909; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_910; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_911; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_912; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_913; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_914; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_915; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_916; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_917; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_918; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_919; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_920; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_921; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_922; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_923; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_924; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_925; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_926; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_927; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_928; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_929; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_930; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_931; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_932; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_933; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_934; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_935; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_936; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_937; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_938; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_939; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_940; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_941; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_942; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_943; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_944; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_945; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_946; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_947; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_948; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_949; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_950; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_951; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_952; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_953; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_954; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_955; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_956; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_957; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_958; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_959; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_960; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_961; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_962; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_963; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_964; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_965; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_966; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_967; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_968; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_969; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_970; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_971; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_972; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_973; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_974; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_975; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_976; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_977; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_978; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_979; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_980; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_981; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_982; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_983; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_984; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_985; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_986; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_987; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_988; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_989; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_990; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_991; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_992; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_993; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_994; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_995; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_996; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_997; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_998; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_999; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1000; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1001; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1002; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1003; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1004; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1005; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1006; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1007; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1008; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1009; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1010; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1011; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1012; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1013; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1014; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1015; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1016; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1017; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1018; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1019; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1020; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1021; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1022; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1023; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1024; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1025; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  wire  _GEN_1026; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  reg  wt_actv_vld_0; // @[NV_NVDLA_CMAC_CORE_active.scala 134:30]
  reg [31:0] _RAND_774;
  reg  wt_actv_pvld_out_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_775;
  reg  wt_actv_pvld_out_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_776;
  reg  wt_actv_pvld_out_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_777;
  reg  wt_actv_pvld_out_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_778;
  reg  wt_actv_pvld_out_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_779;
  reg  wt_actv_pvld_out_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_780;
  reg  wt_actv_pvld_out_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_781;
  reg  wt_actv_pvld_out_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_782;
  reg  wt_actv_pvld_out_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_783;
  reg  wt_actv_pvld_out_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_784;
  reg  wt_actv_pvld_out_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_785;
  reg  wt_actv_pvld_out_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_786;
  reg  wt_actv_pvld_out_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_787;
  reg  wt_actv_pvld_out_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_788;
  reg  wt_actv_pvld_out_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_789;
  reg  wt_actv_pvld_out_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_790;
  reg  wt_actv_pvld_out_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_791;
  reg  wt_actv_pvld_out_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_792;
  reg  wt_actv_pvld_out_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_793;
  reg  wt_actv_pvld_out_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_794;
  reg  wt_actv_pvld_out_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_795;
  reg  wt_actv_pvld_out_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_796;
  reg  wt_actv_pvld_out_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_797;
  reg  wt_actv_pvld_out_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_798;
  reg  wt_actv_pvld_out_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_799;
  reg  wt_actv_pvld_out_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_800;
  reg  wt_actv_pvld_out_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_801;
  reg  wt_actv_pvld_out_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_802;
  reg  wt_actv_pvld_out_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_803;
  reg  wt_actv_pvld_out_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_804;
  reg  wt_actv_pvld_out_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_805;
  reg  wt_actv_pvld_out_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_806;
  reg  wt_actv_pvld_out_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_807;
  reg  wt_actv_pvld_out_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_808;
  reg  wt_actv_pvld_out_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_809;
  reg  wt_actv_pvld_out_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_810;
  reg  wt_actv_pvld_out_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_811;
  reg  wt_actv_pvld_out_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_812;
  reg  wt_actv_pvld_out_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_813;
  reg  wt_actv_pvld_out_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_814;
  reg  wt_actv_pvld_out_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_815;
  reg  wt_actv_pvld_out_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_816;
  reg  wt_actv_pvld_out_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_817;
  reg  wt_actv_pvld_out_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_818;
  reg  wt_actv_pvld_out_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_819;
  reg  wt_actv_pvld_out_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_820;
  reg  wt_actv_pvld_out_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_821;
  reg  wt_actv_pvld_out_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_822;
  reg  wt_actv_pvld_out_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_823;
  reg  wt_actv_pvld_out_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_824;
  reg  wt_actv_pvld_out_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_825;
  reg  wt_actv_pvld_out_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_826;
  reg  wt_actv_pvld_out_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_827;
  reg  wt_actv_pvld_out_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_828;
  reg  wt_actv_pvld_out_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_829;
  reg  wt_actv_pvld_out_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_830;
  reg  wt_actv_pvld_out_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_831;
  reg  wt_actv_pvld_out_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_832;
  reg  wt_actv_pvld_out_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_833;
  reg  wt_actv_pvld_out_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_834;
  reg  wt_actv_pvld_out_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_835;
  reg  wt_actv_pvld_out_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_836;
  reg  wt_actv_pvld_out_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_837;
  reg  wt_actv_pvld_out_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_838;
  reg  wt_actv_pvld_out_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_839;
  reg  wt_actv_pvld_out_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_840;
  reg  wt_actv_pvld_out_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_841;
  reg  wt_actv_pvld_out_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_842;
  reg  wt_actv_pvld_out_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_843;
  reg  wt_actv_pvld_out_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_844;
  reg  wt_actv_pvld_out_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_845;
  reg  wt_actv_pvld_out_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_846;
  reg  wt_actv_pvld_out_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_847;
  reg  wt_actv_pvld_out_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_848;
  reg  wt_actv_pvld_out_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_849;
  reg  wt_actv_pvld_out_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_850;
  reg  wt_actv_pvld_out_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_851;
  reg  wt_actv_pvld_out_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_852;
  reg  wt_actv_pvld_out_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_853;
  reg  wt_actv_pvld_out_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_854;
  reg  wt_actv_pvld_out_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_855;
  reg  wt_actv_pvld_out_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_856;
  reg  wt_actv_pvld_out_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_857;
  reg  wt_actv_pvld_out_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_858;
  reg  wt_actv_pvld_out_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_859;
  reg  wt_actv_pvld_out_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_860;
  reg  wt_actv_pvld_out_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_861;
  reg  wt_actv_pvld_out_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_862;
  reg  wt_actv_pvld_out_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_863;
  reg  wt_actv_pvld_out_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_864;
  reg  wt_actv_pvld_out_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_865;
  reg  wt_actv_pvld_out_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_866;
  reg  wt_actv_pvld_out_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_867;
  reg  wt_actv_pvld_out_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_868;
  reg  wt_actv_pvld_out_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_869;
  reg  wt_actv_pvld_out_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_870;
  reg  wt_actv_pvld_out_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_871;
  reg  wt_actv_pvld_out_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_872;
  reg  wt_actv_pvld_out_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_873;
  reg  wt_actv_pvld_out_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_874;
  reg  wt_actv_pvld_out_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_875;
  reg  wt_actv_pvld_out_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_876;
  reg  wt_actv_pvld_out_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_877;
  reg  wt_actv_pvld_out_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_878;
  reg  wt_actv_pvld_out_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_879;
  reg  wt_actv_pvld_out_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_880;
  reg  wt_actv_pvld_out_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_881;
  reg  wt_actv_pvld_out_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_882;
  reg  wt_actv_pvld_out_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_883;
  reg  wt_actv_pvld_out_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_884;
  reg  wt_actv_pvld_out_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_885;
  reg  wt_actv_pvld_out_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_886;
  reg  wt_actv_pvld_out_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_887;
  reg  wt_actv_pvld_out_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_888;
  reg  wt_actv_pvld_out_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_889;
  reg  wt_actv_pvld_out_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_890;
  reg  wt_actv_pvld_out_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_891;
  reg  wt_actv_pvld_out_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_892;
  reg  wt_actv_pvld_out_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_893;
  reg  wt_actv_pvld_out_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_894;
  reg  wt_actv_pvld_out_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_895;
  reg  wt_actv_pvld_out_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_896;
  reg  wt_actv_pvld_out_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_897;
  reg  wt_actv_pvld_out_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_898;
  reg  wt_actv_pvld_out_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_899;
  reg  wt_actv_pvld_out_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_900;
  reg  wt_actv_pvld_out_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_901;
  reg  wt_actv_pvld_out_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 135:35]
  reg [31:0] _RAND_902;
  reg  wt_actv_nz_out_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_903;
  reg  wt_actv_nz_out_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_904;
  reg  wt_actv_nz_out_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_905;
  reg  wt_actv_nz_out_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_906;
  reg  wt_actv_nz_out_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_907;
  reg  wt_actv_nz_out_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_908;
  reg  wt_actv_nz_out_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_909;
  reg  wt_actv_nz_out_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_910;
  reg  wt_actv_nz_out_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_911;
  reg  wt_actv_nz_out_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_912;
  reg  wt_actv_nz_out_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_913;
  reg  wt_actv_nz_out_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_914;
  reg  wt_actv_nz_out_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_915;
  reg  wt_actv_nz_out_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_916;
  reg  wt_actv_nz_out_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_917;
  reg  wt_actv_nz_out_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_918;
  reg  wt_actv_nz_out_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_919;
  reg  wt_actv_nz_out_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_920;
  reg  wt_actv_nz_out_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_921;
  reg  wt_actv_nz_out_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_922;
  reg  wt_actv_nz_out_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_923;
  reg  wt_actv_nz_out_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_924;
  reg  wt_actv_nz_out_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_925;
  reg  wt_actv_nz_out_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_926;
  reg  wt_actv_nz_out_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_927;
  reg  wt_actv_nz_out_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_928;
  reg  wt_actv_nz_out_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_929;
  reg  wt_actv_nz_out_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_930;
  reg  wt_actv_nz_out_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_931;
  reg  wt_actv_nz_out_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_932;
  reg  wt_actv_nz_out_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_933;
  reg  wt_actv_nz_out_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_934;
  reg  wt_actv_nz_out_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_935;
  reg  wt_actv_nz_out_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_936;
  reg  wt_actv_nz_out_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_937;
  reg  wt_actv_nz_out_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_938;
  reg  wt_actv_nz_out_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_939;
  reg  wt_actv_nz_out_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_940;
  reg  wt_actv_nz_out_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_941;
  reg  wt_actv_nz_out_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_942;
  reg  wt_actv_nz_out_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_943;
  reg  wt_actv_nz_out_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_944;
  reg  wt_actv_nz_out_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_945;
  reg  wt_actv_nz_out_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_946;
  reg  wt_actv_nz_out_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_947;
  reg  wt_actv_nz_out_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_948;
  reg  wt_actv_nz_out_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_949;
  reg  wt_actv_nz_out_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_950;
  reg  wt_actv_nz_out_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_951;
  reg  wt_actv_nz_out_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_952;
  reg  wt_actv_nz_out_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_953;
  reg  wt_actv_nz_out_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_954;
  reg  wt_actv_nz_out_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_955;
  reg  wt_actv_nz_out_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_956;
  reg  wt_actv_nz_out_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_957;
  reg  wt_actv_nz_out_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_958;
  reg  wt_actv_nz_out_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_959;
  reg  wt_actv_nz_out_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_960;
  reg  wt_actv_nz_out_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_961;
  reg  wt_actv_nz_out_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_962;
  reg  wt_actv_nz_out_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_963;
  reg  wt_actv_nz_out_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_964;
  reg  wt_actv_nz_out_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_965;
  reg  wt_actv_nz_out_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_966;
  reg  wt_actv_nz_out_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_967;
  reg  wt_actv_nz_out_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_968;
  reg  wt_actv_nz_out_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_969;
  reg  wt_actv_nz_out_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_970;
  reg  wt_actv_nz_out_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_971;
  reg  wt_actv_nz_out_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_972;
  reg  wt_actv_nz_out_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_973;
  reg  wt_actv_nz_out_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_974;
  reg  wt_actv_nz_out_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_975;
  reg  wt_actv_nz_out_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_976;
  reg  wt_actv_nz_out_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_977;
  reg  wt_actv_nz_out_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_978;
  reg  wt_actv_nz_out_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_979;
  reg  wt_actv_nz_out_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_980;
  reg  wt_actv_nz_out_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_981;
  reg  wt_actv_nz_out_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_982;
  reg  wt_actv_nz_out_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_983;
  reg  wt_actv_nz_out_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_984;
  reg  wt_actv_nz_out_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_985;
  reg  wt_actv_nz_out_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_986;
  reg  wt_actv_nz_out_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_987;
  reg  wt_actv_nz_out_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_988;
  reg  wt_actv_nz_out_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_989;
  reg  wt_actv_nz_out_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_990;
  reg  wt_actv_nz_out_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_991;
  reg  wt_actv_nz_out_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_992;
  reg  wt_actv_nz_out_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_993;
  reg  wt_actv_nz_out_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_994;
  reg  wt_actv_nz_out_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_995;
  reg  wt_actv_nz_out_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_996;
  reg  wt_actv_nz_out_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_997;
  reg  wt_actv_nz_out_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_998;
  reg  wt_actv_nz_out_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_999;
  reg  wt_actv_nz_out_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1000;
  reg  wt_actv_nz_out_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1001;
  reg  wt_actv_nz_out_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1002;
  reg  wt_actv_nz_out_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1003;
  reg  wt_actv_nz_out_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1004;
  reg  wt_actv_nz_out_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1005;
  reg  wt_actv_nz_out_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1006;
  reg  wt_actv_nz_out_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1007;
  reg  wt_actv_nz_out_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1008;
  reg  wt_actv_nz_out_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1009;
  reg  wt_actv_nz_out_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1010;
  reg  wt_actv_nz_out_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1011;
  reg  wt_actv_nz_out_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1012;
  reg  wt_actv_nz_out_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1013;
  reg  wt_actv_nz_out_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1014;
  reg  wt_actv_nz_out_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1015;
  reg  wt_actv_nz_out_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1016;
  reg  wt_actv_nz_out_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1017;
  reg  wt_actv_nz_out_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1018;
  reg  wt_actv_nz_out_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1019;
  reg  wt_actv_nz_out_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1020;
  reg  wt_actv_nz_out_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1021;
  reg  wt_actv_nz_out_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1022;
  reg  wt_actv_nz_out_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1023;
  reg  wt_actv_nz_out_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1024;
  reg  wt_actv_nz_out_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1025;
  reg  wt_actv_nz_out_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1026;
  reg  wt_actv_nz_out_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1027;
  reg  wt_actv_nz_out_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1028;
  reg  wt_actv_nz_out_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1029;
  reg  wt_actv_nz_out_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 137:33]
  reg [31:0] _RAND_1030;
  reg [7:0] wt_actv_data_out_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1031;
  reg [7:0] wt_actv_data_out_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1032;
  reg [7:0] wt_actv_data_out_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1033;
  reg [7:0] wt_actv_data_out_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1034;
  reg [7:0] wt_actv_data_out_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1035;
  reg [7:0] wt_actv_data_out_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1036;
  reg [7:0] wt_actv_data_out_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1037;
  reg [7:0] wt_actv_data_out_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1038;
  reg [7:0] wt_actv_data_out_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1039;
  reg [7:0] wt_actv_data_out_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1040;
  reg [7:0] wt_actv_data_out_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1041;
  reg [7:0] wt_actv_data_out_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1042;
  reg [7:0] wt_actv_data_out_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1043;
  reg [7:0] wt_actv_data_out_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1044;
  reg [7:0] wt_actv_data_out_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1045;
  reg [7:0] wt_actv_data_out_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1046;
  reg [7:0] wt_actv_data_out_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1047;
  reg [7:0] wt_actv_data_out_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1048;
  reg [7:0] wt_actv_data_out_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1049;
  reg [7:0] wt_actv_data_out_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1050;
  reg [7:0] wt_actv_data_out_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1051;
  reg [7:0] wt_actv_data_out_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1052;
  reg [7:0] wt_actv_data_out_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1053;
  reg [7:0] wt_actv_data_out_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1054;
  reg [7:0] wt_actv_data_out_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1055;
  reg [7:0] wt_actv_data_out_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1056;
  reg [7:0] wt_actv_data_out_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1057;
  reg [7:0] wt_actv_data_out_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1058;
  reg [7:0] wt_actv_data_out_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1059;
  reg [7:0] wt_actv_data_out_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1060;
  reg [7:0] wt_actv_data_out_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1061;
  reg [7:0] wt_actv_data_out_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1062;
  reg [7:0] wt_actv_data_out_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1063;
  reg [7:0] wt_actv_data_out_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1064;
  reg [7:0] wt_actv_data_out_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1065;
  reg [7:0] wt_actv_data_out_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1066;
  reg [7:0] wt_actv_data_out_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1067;
  reg [7:0] wt_actv_data_out_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1068;
  reg [7:0] wt_actv_data_out_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1069;
  reg [7:0] wt_actv_data_out_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1070;
  reg [7:0] wt_actv_data_out_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1071;
  reg [7:0] wt_actv_data_out_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1072;
  reg [7:0] wt_actv_data_out_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1073;
  reg [7:0] wt_actv_data_out_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1074;
  reg [7:0] wt_actv_data_out_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1075;
  reg [7:0] wt_actv_data_out_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1076;
  reg [7:0] wt_actv_data_out_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1077;
  reg [7:0] wt_actv_data_out_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1078;
  reg [7:0] wt_actv_data_out_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1079;
  reg [7:0] wt_actv_data_out_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1080;
  reg [7:0] wt_actv_data_out_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1081;
  reg [7:0] wt_actv_data_out_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1082;
  reg [7:0] wt_actv_data_out_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1083;
  reg [7:0] wt_actv_data_out_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1084;
  reg [7:0] wt_actv_data_out_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1085;
  reg [7:0] wt_actv_data_out_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1086;
  reg [7:0] wt_actv_data_out_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1087;
  reg [7:0] wt_actv_data_out_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1088;
  reg [7:0] wt_actv_data_out_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1089;
  reg [7:0] wt_actv_data_out_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1090;
  reg [7:0] wt_actv_data_out_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1091;
  reg [7:0] wt_actv_data_out_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1092;
  reg [7:0] wt_actv_data_out_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1093;
  reg [7:0] wt_actv_data_out_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1094;
  reg [7:0] wt_actv_data_out_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1095;
  reg [7:0] wt_actv_data_out_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1096;
  reg [7:0] wt_actv_data_out_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1097;
  reg [7:0] wt_actv_data_out_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1098;
  reg [7:0] wt_actv_data_out_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1099;
  reg [7:0] wt_actv_data_out_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1100;
  reg [7:0] wt_actv_data_out_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1101;
  reg [7:0] wt_actv_data_out_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1102;
  reg [7:0] wt_actv_data_out_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1103;
  reg [7:0] wt_actv_data_out_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1104;
  reg [7:0] wt_actv_data_out_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1105;
  reg [7:0] wt_actv_data_out_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1106;
  reg [7:0] wt_actv_data_out_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1107;
  reg [7:0] wt_actv_data_out_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1108;
  reg [7:0] wt_actv_data_out_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1109;
  reg [7:0] wt_actv_data_out_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1110;
  reg [7:0] wt_actv_data_out_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1111;
  reg [7:0] wt_actv_data_out_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1112;
  reg [7:0] wt_actv_data_out_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1113;
  reg [7:0] wt_actv_data_out_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1114;
  reg [7:0] wt_actv_data_out_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1115;
  reg [7:0] wt_actv_data_out_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1116;
  reg [7:0] wt_actv_data_out_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1117;
  reg [7:0] wt_actv_data_out_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1118;
  reg [7:0] wt_actv_data_out_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1119;
  reg [7:0] wt_actv_data_out_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1120;
  reg [7:0] wt_actv_data_out_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1121;
  reg [7:0] wt_actv_data_out_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1122;
  reg [7:0] wt_actv_data_out_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1123;
  reg [7:0] wt_actv_data_out_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1124;
  reg [7:0] wt_actv_data_out_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1125;
  reg [7:0] wt_actv_data_out_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1126;
  reg [7:0] wt_actv_data_out_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1127;
  reg [7:0] wt_actv_data_out_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1128;
  reg [7:0] wt_actv_data_out_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1129;
  reg [7:0] wt_actv_data_out_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1130;
  reg [7:0] wt_actv_data_out_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1131;
  reg [7:0] wt_actv_data_out_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1132;
  reg [7:0] wt_actv_data_out_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1133;
  reg [7:0] wt_actv_data_out_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1134;
  reg [7:0] wt_actv_data_out_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1135;
  reg [7:0] wt_actv_data_out_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1136;
  reg [7:0] wt_actv_data_out_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1137;
  reg [7:0] wt_actv_data_out_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1138;
  reg [7:0] wt_actv_data_out_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1139;
  reg [7:0] wt_actv_data_out_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1140;
  reg [7:0] wt_actv_data_out_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1141;
  reg [7:0] wt_actv_data_out_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1142;
  reg [7:0] wt_actv_data_out_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1143;
  reg [7:0] wt_actv_data_out_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1144;
  reg [7:0] wt_actv_data_out_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1145;
  reg [7:0] wt_actv_data_out_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1146;
  reg [7:0] wt_actv_data_out_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1147;
  reg [7:0] wt_actv_data_out_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1148;
  reg [7:0] wt_actv_data_out_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1149;
  reg [7:0] wt_actv_data_out_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1150;
  reg [7:0] wt_actv_data_out_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1151;
  reg [7:0] wt_actv_data_out_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1152;
  reg [7:0] wt_actv_data_out_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1153;
  reg [7:0] wt_actv_data_out_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1154;
  reg [7:0] wt_actv_data_out_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1155;
  reg [7:0] wt_actv_data_out_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1156;
  reg [7:0] wt_actv_data_out_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1157;
  reg [7:0] wt_actv_data_out_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 138:31]
  reg [31:0] _RAND_1158;
  wire  _T_50631; // @[NV_NVDLA_CMAC_CORE_active.scala 141:78]
  wire  wt_actv_pvld_w_0; // @[NV_NVDLA_CMAC_CORE_active.scala 141:33]
  wire  _T_50633; // @[NV_NVDLA_CMAC_CORE_active.scala 145:42]
  wire [7:0] _GEN_1155; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1156; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1158; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1159; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1161; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1162; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1164; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1165; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1167; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1168; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1170; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1171; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1173; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1174; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1176; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1177; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1179; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1180; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1182; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1183; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1185; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1186; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1188; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1189; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1191; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1192; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1194; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1195; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1197; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1198; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1200; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1201; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1203; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1204; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1206; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1207; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1209; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1210; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1212; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1213; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1215; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1216; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1218; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1219; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1221; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1222; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1224; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1225; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1227; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1228; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1230; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1231; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1233; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1234; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1236; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1237; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1239; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1240; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1242; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1243; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1245; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1246; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1248; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1249; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1251; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1252; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1254; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1255; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1257; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1258; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1260; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1261; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1263; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1264; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1266; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1267; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1269; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1270; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1272; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1273; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1275; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1276; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1278; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1279; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1281; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1282; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1284; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1285; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1287; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1288; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1290; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1291; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1293; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1294; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1296; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1297; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1299; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1300; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1302; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1303; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1305; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1306; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1308; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1309; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1311; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1312; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1314; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1315; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1317; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1318; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1320; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1321; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1323; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1324; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1326; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1327; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1329; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1330; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1332; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1333; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1335; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1336; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1338; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1339; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1341; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1342; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1344; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1345; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1347; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1348; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1350; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1351; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1353; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1354; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1356; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1357; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1359; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1360; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1362; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1363; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1365; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1366; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1368; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1369; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1371; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1372; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1374; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1375; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1377; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1378; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1380; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1381; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1383; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1384; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1386; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1387; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1389; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1390; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1392; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1393; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1395; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1396; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1398; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1399; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1401; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1402; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1404; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1405; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1407; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1408; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1410; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1411; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1413; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1414; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1416; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1417; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1419; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1420; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1422; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1423; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1425; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1426; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1428; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1429; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1431; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1432; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1434; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1435; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1437; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1438; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1440; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1441; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1443; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1444; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1446; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1447; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1449; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1450; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1452; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1453; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1455; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1456; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1458; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1459; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1461; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1462; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1464; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1465; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1467; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1468; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1470; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1471; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1473; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1474; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1476; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1477; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1479; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1480; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1482; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1483; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1485; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1486; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1488; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1489; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1491; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1492; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1494; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1495; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1497; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1498; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1500; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1501; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1503; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1504; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1506; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1507; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1509; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1510; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1512; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1513; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1515; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1516; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1518; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1519; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1521; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1522; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1524; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1525; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1527; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1528; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1530; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1531; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1533; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1534; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  wire [7:0] _GEN_1536; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  wire  _GEN_1537; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  reg [7:0] dat_actv_data_reg_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1159;
  reg [7:0] dat_actv_data_reg_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1160;
  reg [7:0] dat_actv_data_reg_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1161;
  reg [7:0] dat_actv_data_reg_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1162;
  reg [7:0] dat_actv_data_reg_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1163;
  reg [7:0] dat_actv_data_reg_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1164;
  reg [7:0] dat_actv_data_reg_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1165;
  reg [7:0] dat_actv_data_reg_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1166;
  reg [7:0] dat_actv_data_reg_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1167;
  reg [7:0] dat_actv_data_reg_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1168;
  reg [7:0] dat_actv_data_reg_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1169;
  reg [7:0] dat_actv_data_reg_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1170;
  reg [7:0] dat_actv_data_reg_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1171;
  reg [7:0] dat_actv_data_reg_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1172;
  reg [7:0] dat_actv_data_reg_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1173;
  reg [7:0] dat_actv_data_reg_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1174;
  reg [7:0] dat_actv_data_reg_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1175;
  reg [7:0] dat_actv_data_reg_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1176;
  reg [7:0] dat_actv_data_reg_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1177;
  reg [7:0] dat_actv_data_reg_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1178;
  reg [7:0] dat_actv_data_reg_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1179;
  reg [7:0] dat_actv_data_reg_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1180;
  reg [7:0] dat_actv_data_reg_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1181;
  reg [7:0] dat_actv_data_reg_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1182;
  reg [7:0] dat_actv_data_reg_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1183;
  reg [7:0] dat_actv_data_reg_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1184;
  reg [7:0] dat_actv_data_reg_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1185;
  reg [7:0] dat_actv_data_reg_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1186;
  reg [7:0] dat_actv_data_reg_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1187;
  reg [7:0] dat_actv_data_reg_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1188;
  reg [7:0] dat_actv_data_reg_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1189;
  reg [7:0] dat_actv_data_reg_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1190;
  reg [7:0] dat_actv_data_reg_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1191;
  reg [7:0] dat_actv_data_reg_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1192;
  reg [7:0] dat_actv_data_reg_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1193;
  reg [7:0] dat_actv_data_reg_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1194;
  reg [7:0] dat_actv_data_reg_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1195;
  reg [7:0] dat_actv_data_reg_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1196;
  reg [7:0] dat_actv_data_reg_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1197;
  reg [7:0] dat_actv_data_reg_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1198;
  reg [7:0] dat_actv_data_reg_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1199;
  reg [7:0] dat_actv_data_reg_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1200;
  reg [7:0] dat_actv_data_reg_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1201;
  reg [7:0] dat_actv_data_reg_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1202;
  reg [7:0] dat_actv_data_reg_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1203;
  reg [7:0] dat_actv_data_reg_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1204;
  reg [7:0] dat_actv_data_reg_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1205;
  reg [7:0] dat_actv_data_reg_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1206;
  reg [7:0] dat_actv_data_reg_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1207;
  reg [7:0] dat_actv_data_reg_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1208;
  reg [7:0] dat_actv_data_reg_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1209;
  reg [7:0] dat_actv_data_reg_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1210;
  reg [7:0] dat_actv_data_reg_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1211;
  reg [7:0] dat_actv_data_reg_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1212;
  reg [7:0] dat_actv_data_reg_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1213;
  reg [7:0] dat_actv_data_reg_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1214;
  reg [7:0] dat_actv_data_reg_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1215;
  reg [7:0] dat_actv_data_reg_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1216;
  reg [7:0] dat_actv_data_reg_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1217;
  reg [7:0] dat_actv_data_reg_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1218;
  reg [7:0] dat_actv_data_reg_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1219;
  reg [7:0] dat_actv_data_reg_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1220;
  reg [7:0] dat_actv_data_reg_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1221;
  reg [7:0] dat_actv_data_reg_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1222;
  reg [7:0] dat_actv_data_reg_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1223;
  reg [7:0] dat_actv_data_reg_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1224;
  reg [7:0] dat_actv_data_reg_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1225;
  reg [7:0] dat_actv_data_reg_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1226;
  reg [7:0] dat_actv_data_reg_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1227;
  reg [7:0] dat_actv_data_reg_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1228;
  reg [7:0] dat_actv_data_reg_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1229;
  reg [7:0] dat_actv_data_reg_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1230;
  reg [7:0] dat_actv_data_reg_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1231;
  reg [7:0] dat_actv_data_reg_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1232;
  reg [7:0] dat_actv_data_reg_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1233;
  reg [7:0] dat_actv_data_reg_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1234;
  reg [7:0] dat_actv_data_reg_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1235;
  reg [7:0] dat_actv_data_reg_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1236;
  reg [7:0] dat_actv_data_reg_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1237;
  reg [7:0] dat_actv_data_reg_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1238;
  reg [7:0] dat_actv_data_reg_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1239;
  reg [7:0] dat_actv_data_reg_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1240;
  reg [7:0] dat_actv_data_reg_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1241;
  reg [7:0] dat_actv_data_reg_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1242;
  reg [7:0] dat_actv_data_reg_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1243;
  reg [7:0] dat_actv_data_reg_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1244;
  reg [7:0] dat_actv_data_reg_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1245;
  reg [7:0] dat_actv_data_reg_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1246;
  reg [7:0] dat_actv_data_reg_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1247;
  reg [7:0] dat_actv_data_reg_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1248;
  reg [7:0] dat_actv_data_reg_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1249;
  reg [7:0] dat_actv_data_reg_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1250;
  reg [7:0] dat_actv_data_reg_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1251;
  reg [7:0] dat_actv_data_reg_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1252;
  reg [7:0] dat_actv_data_reg_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1253;
  reg [7:0] dat_actv_data_reg_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1254;
  reg [7:0] dat_actv_data_reg_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1255;
  reg [7:0] dat_actv_data_reg_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1256;
  reg [7:0] dat_actv_data_reg_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1257;
  reg [7:0] dat_actv_data_reg_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1258;
  reg [7:0] dat_actv_data_reg_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1259;
  reg [7:0] dat_actv_data_reg_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1260;
  reg [7:0] dat_actv_data_reg_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1261;
  reg [7:0] dat_actv_data_reg_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1262;
  reg [7:0] dat_actv_data_reg_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1263;
  reg [7:0] dat_actv_data_reg_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1264;
  reg [7:0] dat_actv_data_reg_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1265;
  reg [7:0] dat_actv_data_reg_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1266;
  reg [7:0] dat_actv_data_reg_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1267;
  reg [7:0] dat_actv_data_reg_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1268;
  reg [7:0] dat_actv_data_reg_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1269;
  reg [7:0] dat_actv_data_reg_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1270;
  reg [7:0] dat_actv_data_reg_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1271;
  reg [7:0] dat_actv_data_reg_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1272;
  reg [7:0] dat_actv_data_reg_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1273;
  reg [7:0] dat_actv_data_reg_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1274;
  reg [7:0] dat_actv_data_reg_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1275;
  reg [7:0] dat_actv_data_reg_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1276;
  reg [7:0] dat_actv_data_reg_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1277;
  reg [7:0] dat_actv_data_reg_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1278;
  reg [7:0] dat_actv_data_reg_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1279;
  reg [7:0] dat_actv_data_reg_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1280;
  reg [7:0] dat_actv_data_reg_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1281;
  reg [7:0] dat_actv_data_reg_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1282;
  reg [7:0] dat_actv_data_reg_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1283;
  reg [7:0] dat_actv_data_reg_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1284;
  reg [7:0] dat_actv_data_reg_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1285;
  reg [7:0] dat_actv_data_reg_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 159:32]
  reg [31:0] _RAND_1286;
  reg  dat_actv_nz_reg_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1287;
  reg  dat_actv_nz_reg_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1288;
  reg  dat_actv_nz_reg_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1289;
  reg  dat_actv_nz_reg_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1290;
  reg  dat_actv_nz_reg_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1291;
  reg  dat_actv_nz_reg_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1292;
  reg  dat_actv_nz_reg_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1293;
  reg  dat_actv_nz_reg_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1294;
  reg  dat_actv_nz_reg_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1295;
  reg  dat_actv_nz_reg_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1296;
  reg  dat_actv_nz_reg_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1297;
  reg  dat_actv_nz_reg_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1298;
  reg  dat_actv_nz_reg_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1299;
  reg  dat_actv_nz_reg_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1300;
  reg  dat_actv_nz_reg_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1301;
  reg  dat_actv_nz_reg_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1302;
  reg  dat_actv_nz_reg_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1303;
  reg  dat_actv_nz_reg_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1304;
  reg  dat_actv_nz_reg_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1305;
  reg  dat_actv_nz_reg_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1306;
  reg  dat_actv_nz_reg_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1307;
  reg  dat_actv_nz_reg_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1308;
  reg  dat_actv_nz_reg_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1309;
  reg  dat_actv_nz_reg_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1310;
  reg  dat_actv_nz_reg_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1311;
  reg  dat_actv_nz_reg_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1312;
  reg  dat_actv_nz_reg_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1313;
  reg  dat_actv_nz_reg_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1314;
  reg  dat_actv_nz_reg_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1315;
  reg  dat_actv_nz_reg_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1316;
  reg  dat_actv_nz_reg_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1317;
  reg  dat_actv_nz_reg_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1318;
  reg  dat_actv_nz_reg_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1319;
  reg  dat_actv_nz_reg_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1320;
  reg  dat_actv_nz_reg_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1321;
  reg  dat_actv_nz_reg_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1322;
  reg  dat_actv_nz_reg_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1323;
  reg  dat_actv_nz_reg_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1324;
  reg  dat_actv_nz_reg_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1325;
  reg  dat_actv_nz_reg_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1326;
  reg  dat_actv_nz_reg_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1327;
  reg  dat_actv_nz_reg_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1328;
  reg  dat_actv_nz_reg_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1329;
  reg  dat_actv_nz_reg_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1330;
  reg  dat_actv_nz_reg_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1331;
  reg  dat_actv_nz_reg_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1332;
  reg  dat_actv_nz_reg_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1333;
  reg  dat_actv_nz_reg_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1334;
  reg  dat_actv_nz_reg_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1335;
  reg  dat_actv_nz_reg_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1336;
  reg  dat_actv_nz_reg_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1337;
  reg  dat_actv_nz_reg_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1338;
  reg  dat_actv_nz_reg_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1339;
  reg  dat_actv_nz_reg_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1340;
  reg  dat_actv_nz_reg_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1341;
  reg  dat_actv_nz_reg_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1342;
  reg  dat_actv_nz_reg_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1343;
  reg  dat_actv_nz_reg_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1344;
  reg  dat_actv_nz_reg_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1345;
  reg  dat_actv_nz_reg_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1346;
  reg  dat_actv_nz_reg_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1347;
  reg  dat_actv_nz_reg_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1348;
  reg  dat_actv_nz_reg_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1349;
  reg  dat_actv_nz_reg_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1350;
  reg  dat_actv_nz_reg_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1351;
  reg  dat_actv_nz_reg_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1352;
  reg  dat_actv_nz_reg_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1353;
  reg  dat_actv_nz_reg_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1354;
  reg  dat_actv_nz_reg_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1355;
  reg  dat_actv_nz_reg_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1356;
  reg  dat_actv_nz_reg_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1357;
  reg  dat_actv_nz_reg_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1358;
  reg  dat_actv_nz_reg_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1359;
  reg  dat_actv_nz_reg_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1360;
  reg  dat_actv_nz_reg_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1361;
  reg  dat_actv_nz_reg_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1362;
  reg  dat_actv_nz_reg_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1363;
  reg  dat_actv_nz_reg_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1364;
  reg  dat_actv_nz_reg_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1365;
  reg  dat_actv_nz_reg_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1366;
  reg  dat_actv_nz_reg_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1367;
  reg  dat_actv_nz_reg_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1368;
  reg  dat_actv_nz_reg_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1369;
  reg  dat_actv_nz_reg_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1370;
  reg  dat_actv_nz_reg_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1371;
  reg  dat_actv_nz_reg_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1372;
  reg  dat_actv_nz_reg_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1373;
  reg  dat_actv_nz_reg_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1374;
  reg  dat_actv_nz_reg_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1375;
  reg  dat_actv_nz_reg_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1376;
  reg  dat_actv_nz_reg_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1377;
  reg  dat_actv_nz_reg_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1378;
  reg  dat_actv_nz_reg_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1379;
  reg  dat_actv_nz_reg_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1380;
  reg  dat_actv_nz_reg_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1381;
  reg  dat_actv_nz_reg_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1382;
  reg  dat_actv_nz_reg_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1383;
  reg  dat_actv_nz_reg_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1384;
  reg  dat_actv_nz_reg_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1385;
  reg  dat_actv_nz_reg_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1386;
  reg  dat_actv_nz_reg_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1387;
  reg  dat_actv_nz_reg_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1388;
  reg  dat_actv_nz_reg_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1389;
  reg  dat_actv_nz_reg_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1390;
  reg  dat_actv_nz_reg_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1391;
  reg  dat_actv_nz_reg_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1392;
  reg  dat_actv_nz_reg_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1393;
  reg  dat_actv_nz_reg_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1394;
  reg  dat_actv_nz_reg_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1395;
  reg  dat_actv_nz_reg_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1396;
  reg  dat_actv_nz_reg_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1397;
  reg  dat_actv_nz_reg_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1398;
  reg  dat_actv_nz_reg_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1399;
  reg  dat_actv_nz_reg_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1400;
  reg  dat_actv_nz_reg_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1401;
  reg  dat_actv_nz_reg_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1402;
  reg  dat_actv_nz_reg_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1403;
  reg  dat_actv_nz_reg_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1404;
  reg  dat_actv_nz_reg_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1405;
  reg  dat_actv_nz_reg_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1406;
  reg  dat_actv_nz_reg_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1407;
  reg  dat_actv_nz_reg_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1408;
  reg  dat_actv_nz_reg_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1409;
  reg  dat_actv_nz_reg_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1410;
  reg  dat_actv_nz_reg_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1411;
  reg  dat_actv_nz_reg_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1412;
  reg  dat_actv_nz_reg_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1413;
  reg  dat_actv_nz_reg_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 160:34]
  reg [31:0] _RAND_1414;
  reg  dat_actv_pvld_reg_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1415;
  reg  dat_actv_pvld_reg_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1416;
  reg  dat_actv_pvld_reg_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1417;
  reg  dat_actv_pvld_reg_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1418;
  reg  dat_actv_pvld_reg_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1419;
  reg  dat_actv_pvld_reg_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1420;
  reg  dat_actv_pvld_reg_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1421;
  reg  dat_actv_pvld_reg_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1422;
  reg  dat_actv_pvld_reg_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1423;
  reg  dat_actv_pvld_reg_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1424;
  reg  dat_actv_pvld_reg_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1425;
  reg  dat_actv_pvld_reg_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1426;
  reg  dat_actv_pvld_reg_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1427;
  reg  dat_actv_pvld_reg_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1428;
  reg  dat_actv_pvld_reg_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1429;
  reg  dat_actv_pvld_reg_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1430;
  reg  dat_actv_pvld_reg_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1431;
  reg  dat_actv_pvld_reg_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1432;
  reg  dat_actv_pvld_reg_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1433;
  reg  dat_actv_pvld_reg_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1434;
  reg  dat_actv_pvld_reg_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1435;
  reg  dat_actv_pvld_reg_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1436;
  reg  dat_actv_pvld_reg_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1437;
  reg  dat_actv_pvld_reg_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1438;
  reg  dat_actv_pvld_reg_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1439;
  reg  dat_actv_pvld_reg_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1440;
  reg  dat_actv_pvld_reg_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1441;
  reg  dat_actv_pvld_reg_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1442;
  reg  dat_actv_pvld_reg_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1443;
  reg  dat_actv_pvld_reg_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1444;
  reg  dat_actv_pvld_reg_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1445;
  reg  dat_actv_pvld_reg_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1446;
  reg  dat_actv_pvld_reg_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1447;
  reg  dat_actv_pvld_reg_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1448;
  reg  dat_actv_pvld_reg_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1449;
  reg  dat_actv_pvld_reg_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1450;
  reg  dat_actv_pvld_reg_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1451;
  reg  dat_actv_pvld_reg_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1452;
  reg  dat_actv_pvld_reg_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1453;
  reg  dat_actv_pvld_reg_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1454;
  reg  dat_actv_pvld_reg_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1455;
  reg  dat_actv_pvld_reg_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1456;
  reg  dat_actv_pvld_reg_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1457;
  reg  dat_actv_pvld_reg_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1458;
  reg  dat_actv_pvld_reg_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1459;
  reg  dat_actv_pvld_reg_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1460;
  reg  dat_actv_pvld_reg_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1461;
  reg  dat_actv_pvld_reg_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1462;
  reg  dat_actv_pvld_reg_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1463;
  reg  dat_actv_pvld_reg_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1464;
  reg  dat_actv_pvld_reg_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1465;
  reg  dat_actv_pvld_reg_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1466;
  reg  dat_actv_pvld_reg_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1467;
  reg  dat_actv_pvld_reg_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1468;
  reg  dat_actv_pvld_reg_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1469;
  reg  dat_actv_pvld_reg_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1470;
  reg  dat_actv_pvld_reg_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1471;
  reg  dat_actv_pvld_reg_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1472;
  reg  dat_actv_pvld_reg_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1473;
  reg  dat_actv_pvld_reg_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1474;
  reg  dat_actv_pvld_reg_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1475;
  reg  dat_actv_pvld_reg_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1476;
  reg  dat_actv_pvld_reg_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1477;
  reg  dat_actv_pvld_reg_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1478;
  reg  dat_actv_pvld_reg_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1479;
  reg  dat_actv_pvld_reg_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1480;
  reg  dat_actv_pvld_reg_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1481;
  reg  dat_actv_pvld_reg_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1482;
  reg  dat_actv_pvld_reg_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1483;
  reg  dat_actv_pvld_reg_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1484;
  reg  dat_actv_pvld_reg_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1485;
  reg  dat_actv_pvld_reg_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1486;
  reg  dat_actv_pvld_reg_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1487;
  reg  dat_actv_pvld_reg_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1488;
  reg  dat_actv_pvld_reg_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1489;
  reg  dat_actv_pvld_reg_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1490;
  reg  dat_actv_pvld_reg_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1491;
  reg  dat_actv_pvld_reg_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1492;
  reg  dat_actv_pvld_reg_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1493;
  reg  dat_actv_pvld_reg_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1494;
  reg  dat_actv_pvld_reg_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1495;
  reg  dat_actv_pvld_reg_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1496;
  reg  dat_actv_pvld_reg_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1497;
  reg  dat_actv_pvld_reg_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1498;
  reg  dat_actv_pvld_reg_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1499;
  reg  dat_actv_pvld_reg_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1500;
  reg  dat_actv_pvld_reg_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1501;
  reg  dat_actv_pvld_reg_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1502;
  reg  dat_actv_pvld_reg_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1503;
  reg  dat_actv_pvld_reg_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1504;
  reg  dat_actv_pvld_reg_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1505;
  reg  dat_actv_pvld_reg_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1506;
  reg  dat_actv_pvld_reg_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1507;
  reg  dat_actv_pvld_reg_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1508;
  reg  dat_actv_pvld_reg_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1509;
  reg  dat_actv_pvld_reg_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1510;
  reg  dat_actv_pvld_reg_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1511;
  reg  dat_actv_pvld_reg_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1512;
  reg  dat_actv_pvld_reg_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1513;
  reg  dat_actv_pvld_reg_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1514;
  reg  dat_actv_pvld_reg_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1515;
  reg  dat_actv_pvld_reg_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1516;
  reg  dat_actv_pvld_reg_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1517;
  reg  dat_actv_pvld_reg_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1518;
  reg  dat_actv_pvld_reg_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1519;
  reg  dat_actv_pvld_reg_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1520;
  reg  dat_actv_pvld_reg_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1521;
  reg  dat_actv_pvld_reg_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1522;
  reg  dat_actv_pvld_reg_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1523;
  reg  dat_actv_pvld_reg_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1524;
  reg  dat_actv_pvld_reg_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1525;
  reg  dat_actv_pvld_reg_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1526;
  reg  dat_actv_pvld_reg_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1527;
  reg  dat_actv_pvld_reg_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1528;
  reg  dat_actv_pvld_reg_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1529;
  reg  dat_actv_pvld_reg_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1530;
  reg  dat_actv_pvld_reg_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1531;
  reg  dat_actv_pvld_reg_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1532;
  reg  dat_actv_pvld_reg_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1533;
  reg  dat_actv_pvld_reg_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1534;
  reg  dat_actv_pvld_reg_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1535;
  reg  dat_actv_pvld_reg_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1536;
  reg  dat_actv_pvld_reg_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1537;
  reg  dat_actv_pvld_reg_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1538;
  reg  dat_actv_pvld_reg_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1539;
  reg  dat_actv_pvld_reg_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1540;
  reg  dat_actv_pvld_reg_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1541;
  reg  dat_actv_pvld_reg_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 161:36]
  reg [31:0] _RAND_1542;
  wire  _GEN_1539; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1540; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1541; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1542; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1543; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1544; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1545; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1546; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1547; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1548; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1549; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1550; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1551; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1552; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1553; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1554; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1555; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1556; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1557; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1558; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1559; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1560; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1561; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1562; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1563; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1564; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1565; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1566; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1567; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1568; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1569; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1570; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1571; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1572; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1573; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1574; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1575; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1576; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1577; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1578; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1579; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1580; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1581; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1582; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1583; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1584; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1585; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1586; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1587; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1588; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1589; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1590; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1591; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1592; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1593; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1594; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1595; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1596; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1597; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1598; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1599; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1600; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1601; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1602; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1603; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1604; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1605; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1606; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1607; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1608; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1609; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1610; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1611; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1612; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1613; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1614; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1615; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1616; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1617; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1618; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1619; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1620; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1621; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1622; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1623; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1624; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1625; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1626; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1627; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1628; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1629; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1630; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1631; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1632; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1633; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1634; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1635; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1636; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1637; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1638; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1639; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1640; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1641; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1642; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1643; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1644; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1645; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1646; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1647; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1648; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1649; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1650; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1651; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1652; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1653; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1654; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1655; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1656; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1657; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1658; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1659; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1660; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1661; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1662; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1663; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1664; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1665; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _GEN_1666; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  wire  _T_73569; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73570; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73571; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73572; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73573; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73574; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73575; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73576; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73577; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73578; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73579; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73580; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73581; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73582; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73583; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73584; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73585; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73586; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73587; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73588; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73589; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73590; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73591; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73592; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73593; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73594; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73595; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73596; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73597; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73598; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73599; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73600; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73601; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73602; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73603; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73604; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73605; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73606; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73607; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73608; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73609; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73610; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73611; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73612; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73613; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73614; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73615; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73616; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73617; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73618; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73619; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73620; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73621; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73622; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73623; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73624; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73625; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73626; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73627; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73628; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73629; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73630; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73631; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73632; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73633; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73634; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73635; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73636; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73637; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73638; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73639; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73640; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73641; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73642; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73643; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73644; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73645; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73646; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73647; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73648; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73649; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73650; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73651; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73652; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73653; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73654; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73655; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73656; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73657; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73658; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73659; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73660; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73661; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73662; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73663; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73664; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73665; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73666; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73667; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73668; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73669; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73670; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73671; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73672; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73673; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73674; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73675; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73676; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73677; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73678; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73679; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73680; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73681; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73682; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73683; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73684; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73685; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73686; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73687; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73688; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73689; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73690; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73691; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73692; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73693; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73694; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73695; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  wire  _T_73696; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _GEN_0 = io_in_wt_mask_0 ? io_in_wt_data_0 : wt_pre_data_0; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_1 = io_in_wt_mask_1 ? io_in_wt_data_1 : wt_pre_data_1; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_2 = io_in_wt_mask_2 ? io_in_wt_data_2 : wt_pre_data_2; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_3 = io_in_wt_mask_3 ? io_in_wt_data_3 : wt_pre_data_3; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_4 = io_in_wt_mask_4 ? io_in_wt_data_4 : wt_pre_data_4; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_5 = io_in_wt_mask_5 ? io_in_wt_data_5 : wt_pre_data_5; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_6 = io_in_wt_mask_6 ? io_in_wt_data_6 : wt_pre_data_6; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_7 = io_in_wt_mask_7 ? io_in_wt_data_7 : wt_pre_data_7; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_8 = io_in_wt_mask_8 ? io_in_wt_data_8 : wt_pre_data_8; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_9 = io_in_wt_mask_9 ? io_in_wt_data_9 : wt_pre_data_9; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_10 = io_in_wt_mask_10 ? io_in_wt_data_10 : wt_pre_data_10; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_11 = io_in_wt_mask_11 ? io_in_wt_data_11 : wt_pre_data_11; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_12 = io_in_wt_mask_12 ? io_in_wt_data_12 : wt_pre_data_12; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_13 = io_in_wt_mask_13 ? io_in_wt_data_13 : wt_pre_data_13; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_14 = io_in_wt_mask_14 ? io_in_wt_data_14 : wt_pre_data_14; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_15 = io_in_wt_mask_15 ? io_in_wt_data_15 : wt_pre_data_15; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_16 = io_in_wt_mask_16 ? io_in_wt_data_16 : wt_pre_data_16; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_17 = io_in_wt_mask_17 ? io_in_wt_data_17 : wt_pre_data_17; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_18 = io_in_wt_mask_18 ? io_in_wt_data_18 : wt_pre_data_18; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_19 = io_in_wt_mask_19 ? io_in_wt_data_19 : wt_pre_data_19; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_20 = io_in_wt_mask_20 ? io_in_wt_data_20 : wt_pre_data_20; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_21 = io_in_wt_mask_21 ? io_in_wt_data_21 : wt_pre_data_21; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_22 = io_in_wt_mask_22 ? io_in_wt_data_22 : wt_pre_data_22; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_23 = io_in_wt_mask_23 ? io_in_wt_data_23 : wt_pre_data_23; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_24 = io_in_wt_mask_24 ? io_in_wt_data_24 : wt_pre_data_24; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_25 = io_in_wt_mask_25 ? io_in_wt_data_25 : wt_pre_data_25; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_26 = io_in_wt_mask_26 ? io_in_wt_data_26 : wt_pre_data_26; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_27 = io_in_wt_mask_27 ? io_in_wt_data_27 : wt_pre_data_27; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_28 = io_in_wt_mask_28 ? io_in_wt_data_28 : wt_pre_data_28; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_29 = io_in_wt_mask_29 ? io_in_wt_data_29 : wt_pre_data_29; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_30 = io_in_wt_mask_30 ? io_in_wt_data_30 : wt_pre_data_30; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_31 = io_in_wt_mask_31 ? io_in_wt_data_31 : wt_pre_data_31; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_32 = io_in_wt_mask_32 ? io_in_wt_data_32 : wt_pre_data_32; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_33 = io_in_wt_mask_33 ? io_in_wt_data_33 : wt_pre_data_33; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_34 = io_in_wt_mask_34 ? io_in_wt_data_34 : wt_pre_data_34; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_35 = io_in_wt_mask_35 ? io_in_wt_data_35 : wt_pre_data_35; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_36 = io_in_wt_mask_36 ? io_in_wt_data_36 : wt_pre_data_36; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_37 = io_in_wt_mask_37 ? io_in_wt_data_37 : wt_pre_data_37; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_38 = io_in_wt_mask_38 ? io_in_wt_data_38 : wt_pre_data_38; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_39 = io_in_wt_mask_39 ? io_in_wt_data_39 : wt_pre_data_39; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_40 = io_in_wt_mask_40 ? io_in_wt_data_40 : wt_pre_data_40; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_41 = io_in_wt_mask_41 ? io_in_wt_data_41 : wt_pre_data_41; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_42 = io_in_wt_mask_42 ? io_in_wt_data_42 : wt_pre_data_42; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_43 = io_in_wt_mask_43 ? io_in_wt_data_43 : wt_pre_data_43; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_44 = io_in_wt_mask_44 ? io_in_wt_data_44 : wt_pre_data_44; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_45 = io_in_wt_mask_45 ? io_in_wt_data_45 : wt_pre_data_45; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_46 = io_in_wt_mask_46 ? io_in_wt_data_46 : wt_pre_data_46; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_47 = io_in_wt_mask_47 ? io_in_wt_data_47 : wt_pre_data_47; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_48 = io_in_wt_mask_48 ? io_in_wt_data_48 : wt_pre_data_48; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_49 = io_in_wt_mask_49 ? io_in_wt_data_49 : wt_pre_data_49; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_50 = io_in_wt_mask_50 ? io_in_wt_data_50 : wt_pre_data_50; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_51 = io_in_wt_mask_51 ? io_in_wt_data_51 : wt_pre_data_51; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_52 = io_in_wt_mask_52 ? io_in_wt_data_52 : wt_pre_data_52; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_53 = io_in_wt_mask_53 ? io_in_wt_data_53 : wt_pre_data_53; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_54 = io_in_wt_mask_54 ? io_in_wt_data_54 : wt_pre_data_54; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_55 = io_in_wt_mask_55 ? io_in_wt_data_55 : wt_pre_data_55; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_56 = io_in_wt_mask_56 ? io_in_wt_data_56 : wt_pre_data_56; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_57 = io_in_wt_mask_57 ? io_in_wt_data_57 : wt_pre_data_57; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_58 = io_in_wt_mask_58 ? io_in_wt_data_58 : wt_pre_data_58; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_59 = io_in_wt_mask_59 ? io_in_wt_data_59 : wt_pre_data_59; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_60 = io_in_wt_mask_60 ? io_in_wt_data_60 : wt_pre_data_60; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_61 = io_in_wt_mask_61 ? io_in_wt_data_61 : wt_pre_data_61; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_62 = io_in_wt_mask_62 ? io_in_wt_data_62 : wt_pre_data_62; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_63 = io_in_wt_mask_63 ? io_in_wt_data_63 : wt_pre_data_63; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_64 = io_in_wt_mask_64 ? io_in_wt_data_64 : wt_pre_data_64; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_65 = io_in_wt_mask_65 ? io_in_wt_data_65 : wt_pre_data_65; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_66 = io_in_wt_mask_66 ? io_in_wt_data_66 : wt_pre_data_66; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_67 = io_in_wt_mask_67 ? io_in_wt_data_67 : wt_pre_data_67; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_68 = io_in_wt_mask_68 ? io_in_wt_data_68 : wt_pre_data_68; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_69 = io_in_wt_mask_69 ? io_in_wt_data_69 : wt_pre_data_69; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_70 = io_in_wt_mask_70 ? io_in_wt_data_70 : wt_pre_data_70; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_71 = io_in_wt_mask_71 ? io_in_wt_data_71 : wt_pre_data_71; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_72 = io_in_wt_mask_72 ? io_in_wt_data_72 : wt_pre_data_72; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_73 = io_in_wt_mask_73 ? io_in_wt_data_73 : wt_pre_data_73; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_74 = io_in_wt_mask_74 ? io_in_wt_data_74 : wt_pre_data_74; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_75 = io_in_wt_mask_75 ? io_in_wt_data_75 : wt_pre_data_75; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_76 = io_in_wt_mask_76 ? io_in_wt_data_76 : wt_pre_data_76; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_77 = io_in_wt_mask_77 ? io_in_wt_data_77 : wt_pre_data_77; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_78 = io_in_wt_mask_78 ? io_in_wt_data_78 : wt_pre_data_78; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_79 = io_in_wt_mask_79 ? io_in_wt_data_79 : wt_pre_data_79; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_80 = io_in_wt_mask_80 ? io_in_wt_data_80 : wt_pre_data_80; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_81 = io_in_wt_mask_81 ? io_in_wt_data_81 : wt_pre_data_81; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_82 = io_in_wt_mask_82 ? io_in_wt_data_82 : wt_pre_data_82; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_83 = io_in_wt_mask_83 ? io_in_wt_data_83 : wt_pre_data_83; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_84 = io_in_wt_mask_84 ? io_in_wt_data_84 : wt_pre_data_84; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_85 = io_in_wt_mask_85 ? io_in_wt_data_85 : wt_pre_data_85; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_86 = io_in_wt_mask_86 ? io_in_wt_data_86 : wt_pre_data_86; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_87 = io_in_wt_mask_87 ? io_in_wt_data_87 : wt_pre_data_87; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_88 = io_in_wt_mask_88 ? io_in_wt_data_88 : wt_pre_data_88; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_89 = io_in_wt_mask_89 ? io_in_wt_data_89 : wt_pre_data_89; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_90 = io_in_wt_mask_90 ? io_in_wt_data_90 : wt_pre_data_90; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_91 = io_in_wt_mask_91 ? io_in_wt_data_91 : wt_pre_data_91; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_92 = io_in_wt_mask_92 ? io_in_wt_data_92 : wt_pre_data_92; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_93 = io_in_wt_mask_93 ? io_in_wt_data_93 : wt_pre_data_93; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_94 = io_in_wt_mask_94 ? io_in_wt_data_94 : wt_pre_data_94; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_95 = io_in_wt_mask_95 ? io_in_wt_data_95 : wt_pre_data_95; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_96 = io_in_wt_mask_96 ? io_in_wt_data_96 : wt_pre_data_96; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_97 = io_in_wt_mask_97 ? io_in_wt_data_97 : wt_pre_data_97; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_98 = io_in_wt_mask_98 ? io_in_wt_data_98 : wt_pre_data_98; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_99 = io_in_wt_mask_99 ? io_in_wt_data_99 : wt_pre_data_99; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_100 = io_in_wt_mask_100 ? io_in_wt_data_100 : wt_pre_data_100; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_101 = io_in_wt_mask_101 ? io_in_wt_data_101 : wt_pre_data_101; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_102 = io_in_wt_mask_102 ? io_in_wt_data_102 : wt_pre_data_102; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_103 = io_in_wt_mask_103 ? io_in_wt_data_103 : wt_pre_data_103; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_104 = io_in_wt_mask_104 ? io_in_wt_data_104 : wt_pre_data_104; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_105 = io_in_wt_mask_105 ? io_in_wt_data_105 : wt_pre_data_105; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_106 = io_in_wt_mask_106 ? io_in_wt_data_106 : wt_pre_data_106; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_107 = io_in_wt_mask_107 ? io_in_wt_data_107 : wt_pre_data_107; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_108 = io_in_wt_mask_108 ? io_in_wt_data_108 : wt_pre_data_108; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_109 = io_in_wt_mask_109 ? io_in_wt_data_109 : wt_pre_data_109; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_110 = io_in_wt_mask_110 ? io_in_wt_data_110 : wt_pre_data_110; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_111 = io_in_wt_mask_111 ? io_in_wt_data_111 : wt_pre_data_111; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_112 = io_in_wt_mask_112 ? io_in_wt_data_112 : wt_pre_data_112; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_113 = io_in_wt_mask_113 ? io_in_wt_data_113 : wt_pre_data_113; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_114 = io_in_wt_mask_114 ? io_in_wt_data_114 : wt_pre_data_114; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_115 = io_in_wt_mask_115 ? io_in_wt_data_115 : wt_pre_data_115; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_116 = io_in_wt_mask_116 ? io_in_wt_data_116 : wt_pre_data_116; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_117 = io_in_wt_mask_117 ? io_in_wt_data_117 : wt_pre_data_117; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_118 = io_in_wt_mask_118 ? io_in_wt_data_118 : wt_pre_data_118; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_119 = io_in_wt_mask_119 ? io_in_wt_data_119 : wt_pre_data_119; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_120 = io_in_wt_mask_120 ? io_in_wt_data_120 : wt_pre_data_120; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_121 = io_in_wt_mask_121 ? io_in_wt_data_121 : wt_pre_data_121; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_122 = io_in_wt_mask_122 ? io_in_wt_data_122 : wt_pre_data_122; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_123 = io_in_wt_mask_123 ? io_in_wt_data_123 : wt_pre_data_123; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_124 = io_in_wt_mask_124 ? io_in_wt_data_124 : wt_pre_data_124; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_125 = io_in_wt_mask_125 ? io_in_wt_data_125 : wt_pre_data_125; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_126 = io_in_wt_mask_126 ? io_in_wt_data_126 : wt_pre_data_126; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_127 = io_in_wt_mask_127 ? io_in_wt_data_127 : wt_pre_data_127; // @[NV_NVDLA_CMAC_CORE_active.scala 75:35]
  assign _GEN_128 = io_in_wt_pvld ? io_in_wt_mask_0 : wt_pre_nz_0; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_129 = io_in_wt_pvld ? io_in_wt_mask_1 : wt_pre_nz_1; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_130 = io_in_wt_pvld ? io_in_wt_mask_2 : wt_pre_nz_2; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_131 = io_in_wt_pvld ? io_in_wt_mask_3 : wt_pre_nz_3; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_132 = io_in_wt_pvld ? io_in_wt_mask_4 : wt_pre_nz_4; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_133 = io_in_wt_pvld ? io_in_wt_mask_5 : wt_pre_nz_5; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_134 = io_in_wt_pvld ? io_in_wt_mask_6 : wt_pre_nz_6; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_135 = io_in_wt_pvld ? io_in_wt_mask_7 : wt_pre_nz_7; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_136 = io_in_wt_pvld ? io_in_wt_mask_8 : wt_pre_nz_8; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_137 = io_in_wt_pvld ? io_in_wt_mask_9 : wt_pre_nz_9; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_138 = io_in_wt_pvld ? io_in_wt_mask_10 : wt_pre_nz_10; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_139 = io_in_wt_pvld ? io_in_wt_mask_11 : wt_pre_nz_11; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_140 = io_in_wt_pvld ? io_in_wt_mask_12 : wt_pre_nz_12; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_141 = io_in_wt_pvld ? io_in_wt_mask_13 : wt_pre_nz_13; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_142 = io_in_wt_pvld ? io_in_wt_mask_14 : wt_pre_nz_14; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_143 = io_in_wt_pvld ? io_in_wt_mask_15 : wt_pre_nz_15; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_144 = io_in_wt_pvld ? io_in_wt_mask_16 : wt_pre_nz_16; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_145 = io_in_wt_pvld ? io_in_wt_mask_17 : wt_pre_nz_17; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_146 = io_in_wt_pvld ? io_in_wt_mask_18 : wt_pre_nz_18; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_147 = io_in_wt_pvld ? io_in_wt_mask_19 : wt_pre_nz_19; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_148 = io_in_wt_pvld ? io_in_wt_mask_20 : wt_pre_nz_20; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_149 = io_in_wt_pvld ? io_in_wt_mask_21 : wt_pre_nz_21; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_150 = io_in_wt_pvld ? io_in_wt_mask_22 : wt_pre_nz_22; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_151 = io_in_wt_pvld ? io_in_wt_mask_23 : wt_pre_nz_23; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_152 = io_in_wt_pvld ? io_in_wt_mask_24 : wt_pre_nz_24; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_153 = io_in_wt_pvld ? io_in_wt_mask_25 : wt_pre_nz_25; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_154 = io_in_wt_pvld ? io_in_wt_mask_26 : wt_pre_nz_26; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_155 = io_in_wt_pvld ? io_in_wt_mask_27 : wt_pre_nz_27; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_156 = io_in_wt_pvld ? io_in_wt_mask_28 : wt_pre_nz_28; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_157 = io_in_wt_pvld ? io_in_wt_mask_29 : wt_pre_nz_29; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_158 = io_in_wt_pvld ? io_in_wt_mask_30 : wt_pre_nz_30; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_159 = io_in_wt_pvld ? io_in_wt_mask_31 : wt_pre_nz_31; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_160 = io_in_wt_pvld ? io_in_wt_mask_32 : wt_pre_nz_32; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_161 = io_in_wt_pvld ? io_in_wt_mask_33 : wt_pre_nz_33; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_162 = io_in_wt_pvld ? io_in_wt_mask_34 : wt_pre_nz_34; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_163 = io_in_wt_pvld ? io_in_wt_mask_35 : wt_pre_nz_35; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_164 = io_in_wt_pvld ? io_in_wt_mask_36 : wt_pre_nz_36; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_165 = io_in_wt_pvld ? io_in_wt_mask_37 : wt_pre_nz_37; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_166 = io_in_wt_pvld ? io_in_wt_mask_38 : wt_pre_nz_38; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_167 = io_in_wt_pvld ? io_in_wt_mask_39 : wt_pre_nz_39; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_168 = io_in_wt_pvld ? io_in_wt_mask_40 : wt_pre_nz_40; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_169 = io_in_wt_pvld ? io_in_wt_mask_41 : wt_pre_nz_41; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_170 = io_in_wt_pvld ? io_in_wt_mask_42 : wt_pre_nz_42; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_171 = io_in_wt_pvld ? io_in_wt_mask_43 : wt_pre_nz_43; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_172 = io_in_wt_pvld ? io_in_wt_mask_44 : wt_pre_nz_44; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_173 = io_in_wt_pvld ? io_in_wt_mask_45 : wt_pre_nz_45; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_174 = io_in_wt_pvld ? io_in_wt_mask_46 : wt_pre_nz_46; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_175 = io_in_wt_pvld ? io_in_wt_mask_47 : wt_pre_nz_47; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_176 = io_in_wt_pvld ? io_in_wt_mask_48 : wt_pre_nz_48; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_177 = io_in_wt_pvld ? io_in_wt_mask_49 : wt_pre_nz_49; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_178 = io_in_wt_pvld ? io_in_wt_mask_50 : wt_pre_nz_50; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_179 = io_in_wt_pvld ? io_in_wt_mask_51 : wt_pre_nz_51; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_180 = io_in_wt_pvld ? io_in_wt_mask_52 : wt_pre_nz_52; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_181 = io_in_wt_pvld ? io_in_wt_mask_53 : wt_pre_nz_53; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_182 = io_in_wt_pvld ? io_in_wt_mask_54 : wt_pre_nz_54; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_183 = io_in_wt_pvld ? io_in_wt_mask_55 : wt_pre_nz_55; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_184 = io_in_wt_pvld ? io_in_wt_mask_56 : wt_pre_nz_56; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_185 = io_in_wt_pvld ? io_in_wt_mask_57 : wt_pre_nz_57; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_186 = io_in_wt_pvld ? io_in_wt_mask_58 : wt_pre_nz_58; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_187 = io_in_wt_pvld ? io_in_wt_mask_59 : wt_pre_nz_59; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_188 = io_in_wt_pvld ? io_in_wt_mask_60 : wt_pre_nz_60; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_189 = io_in_wt_pvld ? io_in_wt_mask_61 : wt_pre_nz_61; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_190 = io_in_wt_pvld ? io_in_wt_mask_62 : wt_pre_nz_62; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_191 = io_in_wt_pvld ? io_in_wt_mask_63 : wt_pre_nz_63; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_192 = io_in_wt_pvld ? io_in_wt_mask_64 : wt_pre_nz_64; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_193 = io_in_wt_pvld ? io_in_wt_mask_65 : wt_pre_nz_65; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_194 = io_in_wt_pvld ? io_in_wt_mask_66 : wt_pre_nz_66; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_195 = io_in_wt_pvld ? io_in_wt_mask_67 : wt_pre_nz_67; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_196 = io_in_wt_pvld ? io_in_wt_mask_68 : wt_pre_nz_68; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_197 = io_in_wt_pvld ? io_in_wt_mask_69 : wt_pre_nz_69; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_198 = io_in_wt_pvld ? io_in_wt_mask_70 : wt_pre_nz_70; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_199 = io_in_wt_pvld ? io_in_wt_mask_71 : wt_pre_nz_71; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_200 = io_in_wt_pvld ? io_in_wt_mask_72 : wt_pre_nz_72; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_201 = io_in_wt_pvld ? io_in_wt_mask_73 : wt_pre_nz_73; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_202 = io_in_wt_pvld ? io_in_wt_mask_74 : wt_pre_nz_74; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_203 = io_in_wt_pvld ? io_in_wt_mask_75 : wt_pre_nz_75; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_204 = io_in_wt_pvld ? io_in_wt_mask_76 : wt_pre_nz_76; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_205 = io_in_wt_pvld ? io_in_wt_mask_77 : wt_pre_nz_77; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_206 = io_in_wt_pvld ? io_in_wt_mask_78 : wt_pre_nz_78; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_207 = io_in_wt_pvld ? io_in_wt_mask_79 : wt_pre_nz_79; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_208 = io_in_wt_pvld ? io_in_wt_mask_80 : wt_pre_nz_80; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_209 = io_in_wt_pvld ? io_in_wt_mask_81 : wt_pre_nz_81; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_210 = io_in_wt_pvld ? io_in_wt_mask_82 : wt_pre_nz_82; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_211 = io_in_wt_pvld ? io_in_wt_mask_83 : wt_pre_nz_83; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_212 = io_in_wt_pvld ? io_in_wt_mask_84 : wt_pre_nz_84; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_213 = io_in_wt_pvld ? io_in_wt_mask_85 : wt_pre_nz_85; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_214 = io_in_wt_pvld ? io_in_wt_mask_86 : wt_pre_nz_86; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_215 = io_in_wt_pvld ? io_in_wt_mask_87 : wt_pre_nz_87; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_216 = io_in_wt_pvld ? io_in_wt_mask_88 : wt_pre_nz_88; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_217 = io_in_wt_pvld ? io_in_wt_mask_89 : wt_pre_nz_89; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_218 = io_in_wt_pvld ? io_in_wt_mask_90 : wt_pre_nz_90; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_219 = io_in_wt_pvld ? io_in_wt_mask_91 : wt_pre_nz_91; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_220 = io_in_wt_pvld ? io_in_wt_mask_92 : wt_pre_nz_92; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_221 = io_in_wt_pvld ? io_in_wt_mask_93 : wt_pre_nz_93; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_222 = io_in_wt_pvld ? io_in_wt_mask_94 : wt_pre_nz_94; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_223 = io_in_wt_pvld ? io_in_wt_mask_95 : wt_pre_nz_95; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_224 = io_in_wt_pvld ? io_in_wt_mask_96 : wt_pre_nz_96; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_225 = io_in_wt_pvld ? io_in_wt_mask_97 : wt_pre_nz_97; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_226 = io_in_wt_pvld ? io_in_wt_mask_98 : wt_pre_nz_98; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_227 = io_in_wt_pvld ? io_in_wt_mask_99 : wt_pre_nz_99; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_228 = io_in_wt_pvld ? io_in_wt_mask_100 : wt_pre_nz_100; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_229 = io_in_wt_pvld ? io_in_wt_mask_101 : wt_pre_nz_101; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_230 = io_in_wt_pvld ? io_in_wt_mask_102 : wt_pre_nz_102; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_231 = io_in_wt_pvld ? io_in_wt_mask_103 : wt_pre_nz_103; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_232 = io_in_wt_pvld ? io_in_wt_mask_104 : wt_pre_nz_104; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_233 = io_in_wt_pvld ? io_in_wt_mask_105 : wt_pre_nz_105; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_234 = io_in_wt_pvld ? io_in_wt_mask_106 : wt_pre_nz_106; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_235 = io_in_wt_pvld ? io_in_wt_mask_107 : wt_pre_nz_107; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_236 = io_in_wt_pvld ? io_in_wt_mask_108 : wt_pre_nz_108; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_237 = io_in_wt_pvld ? io_in_wt_mask_109 : wt_pre_nz_109; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_238 = io_in_wt_pvld ? io_in_wt_mask_110 : wt_pre_nz_110; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_239 = io_in_wt_pvld ? io_in_wt_mask_111 : wt_pre_nz_111; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_240 = io_in_wt_pvld ? io_in_wt_mask_112 : wt_pre_nz_112; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_241 = io_in_wt_pvld ? io_in_wt_mask_113 : wt_pre_nz_113; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_242 = io_in_wt_pvld ? io_in_wt_mask_114 : wt_pre_nz_114; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_243 = io_in_wt_pvld ? io_in_wt_mask_115 : wt_pre_nz_115; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_244 = io_in_wt_pvld ? io_in_wt_mask_116 : wt_pre_nz_116; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_245 = io_in_wt_pvld ? io_in_wt_mask_117 : wt_pre_nz_117; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_246 = io_in_wt_pvld ? io_in_wt_mask_118 : wt_pre_nz_118; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_247 = io_in_wt_pvld ? io_in_wt_mask_119 : wt_pre_nz_119; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_248 = io_in_wt_pvld ? io_in_wt_mask_120 : wt_pre_nz_120; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_249 = io_in_wt_pvld ? io_in_wt_mask_121 : wt_pre_nz_121; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_250 = io_in_wt_pvld ? io_in_wt_mask_122 : wt_pre_nz_122; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_251 = io_in_wt_pvld ? io_in_wt_mask_123 : wt_pre_nz_123; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_252 = io_in_wt_pvld ? io_in_wt_mask_124 : wt_pre_nz_124; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_253 = io_in_wt_pvld ? io_in_wt_mask_125 : wt_pre_nz_125; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_254 = io_in_wt_pvld ? io_in_wt_mask_126 : wt_pre_nz_126; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_255 = io_in_wt_pvld ? io_in_wt_mask_127 : wt_pre_nz_127; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_256 = io_in_wt_pvld ? io_in_wt_sel_0 : wt_pre_sel_0; // @[NV_NVDLA_CMAC_CORE_active.scala 69:24]
  assign _GEN_385 = io_in_dat_mask_0 ? io_in_dat_data_0 : dat_pre_data_0; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_386 = io_in_dat_mask_1 ? io_in_dat_data_1 : dat_pre_data_1; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_387 = io_in_dat_mask_2 ? io_in_dat_data_2 : dat_pre_data_2; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_388 = io_in_dat_mask_3 ? io_in_dat_data_3 : dat_pre_data_3; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_389 = io_in_dat_mask_4 ? io_in_dat_data_4 : dat_pre_data_4; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_390 = io_in_dat_mask_5 ? io_in_dat_data_5 : dat_pre_data_5; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_391 = io_in_dat_mask_6 ? io_in_dat_data_6 : dat_pre_data_6; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_392 = io_in_dat_mask_7 ? io_in_dat_data_7 : dat_pre_data_7; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_393 = io_in_dat_mask_8 ? io_in_dat_data_8 : dat_pre_data_8; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_394 = io_in_dat_mask_9 ? io_in_dat_data_9 : dat_pre_data_9; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_395 = io_in_dat_mask_10 ? io_in_dat_data_10 : dat_pre_data_10; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_396 = io_in_dat_mask_11 ? io_in_dat_data_11 : dat_pre_data_11; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_397 = io_in_dat_mask_12 ? io_in_dat_data_12 : dat_pre_data_12; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_398 = io_in_dat_mask_13 ? io_in_dat_data_13 : dat_pre_data_13; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_399 = io_in_dat_mask_14 ? io_in_dat_data_14 : dat_pre_data_14; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_400 = io_in_dat_mask_15 ? io_in_dat_data_15 : dat_pre_data_15; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_401 = io_in_dat_mask_16 ? io_in_dat_data_16 : dat_pre_data_16; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_402 = io_in_dat_mask_17 ? io_in_dat_data_17 : dat_pre_data_17; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_403 = io_in_dat_mask_18 ? io_in_dat_data_18 : dat_pre_data_18; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_404 = io_in_dat_mask_19 ? io_in_dat_data_19 : dat_pre_data_19; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_405 = io_in_dat_mask_20 ? io_in_dat_data_20 : dat_pre_data_20; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_406 = io_in_dat_mask_21 ? io_in_dat_data_21 : dat_pre_data_21; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_407 = io_in_dat_mask_22 ? io_in_dat_data_22 : dat_pre_data_22; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_408 = io_in_dat_mask_23 ? io_in_dat_data_23 : dat_pre_data_23; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_409 = io_in_dat_mask_24 ? io_in_dat_data_24 : dat_pre_data_24; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_410 = io_in_dat_mask_25 ? io_in_dat_data_25 : dat_pre_data_25; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_411 = io_in_dat_mask_26 ? io_in_dat_data_26 : dat_pre_data_26; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_412 = io_in_dat_mask_27 ? io_in_dat_data_27 : dat_pre_data_27; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_413 = io_in_dat_mask_28 ? io_in_dat_data_28 : dat_pre_data_28; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_414 = io_in_dat_mask_29 ? io_in_dat_data_29 : dat_pre_data_29; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_415 = io_in_dat_mask_30 ? io_in_dat_data_30 : dat_pre_data_30; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_416 = io_in_dat_mask_31 ? io_in_dat_data_31 : dat_pre_data_31; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_417 = io_in_dat_mask_32 ? io_in_dat_data_32 : dat_pre_data_32; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_418 = io_in_dat_mask_33 ? io_in_dat_data_33 : dat_pre_data_33; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_419 = io_in_dat_mask_34 ? io_in_dat_data_34 : dat_pre_data_34; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_420 = io_in_dat_mask_35 ? io_in_dat_data_35 : dat_pre_data_35; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_421 = io_in_dat_mask_36 ? io_in_dat_data_36 : dat_pre_data_36; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_422 = io_in_dat_mask_37 ? io_in_dat_data_37 : dat_pre_data_37; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_423 = io_in_dat_mask_38 ? io_in_dat_data_38 : dat_pre_data_38; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_424 = io_in_dat_mask_39 ? io_in_dat_data_39 : dat_pre_data_39; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_425 = io_in_dat_mask_40 ? io_in_dat_data_40 : dat_pre_data_40; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_426 = io_in_dat_mask_41 ? io_in_dat_data_41 : dat_pre_data_41; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_427 = io_in_dat_mask_42 ? io_in_dat_data_42 : dat_pre_data_42; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_428 = io_in_dat_mask_43 ? io_in_dat_data_43 : dat_pre_data_43; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_429 = io_in_dat_mask_44 ? io_in_dat_data_44 : dat_pre_data_44; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_430 = io_in_dat_mask_45 ? io_in_dat_data_45 : dat_pre_data_45; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_431 = io_in_dat_mask_46 ? io_in_dat_data_46 : dat_pre_data_46; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_432 = io_in_dat_mask_47 ? io_in_dat_data_47 : dat_pre_data_47; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_433 = io_in_dat_mask_48 ? io_in_dat_data_48 : dat_pre_data_48; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_434 = io_in_dat_mask_49 ? io_in_dat_data_49 : dat_pre_data_49; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_435 = io_in_dat_mask_50 ? io_in_dat_data_50 : dat_pre_data_50; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_436 = io_in_dat_mask_51 ? io_in_dat_data_51 : dat_pre_data_51; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_437 = io_in_dat_mask_52 ? io_in_dat_data_52 : dat_pre_data_52; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_438 = io_in_dat_mask_53 ? io_in_dat_data_53 : dat_pre_data_53; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_439 = io_in_dat_mask_54 ? io_in_dat_data_54 : dat_pre_data_54; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_440 = io_in_dat_mask_55 ? io_in_dat_data_55 : dat_pre_data_55; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_441 = io_in_dat_mask_56 ? io_in_dat_data_56 : dat_pre_data_56; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_442 = io_in_dat_mask_57 ? io_in_dat_data_57 : dat_pre_data_57; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_443 = io_in_dat_mask_58 ? io_in_dat_data_58 : dat_pre_data_58; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_444 = io_in_dat_mask_59 ? io_in_dat_data_59 : dat_pre_data_59; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_445 = io_in_dat_mask_60 ? io_in_dat_data_60 : dat_pre_data_60; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_446 = io_in_dat_mask_61 ? io_in_dat_data_61 : dat_pre_data_61; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_447 = io_in_dat_mask_62 ? io_in_dat_data_62 : dat_pre_data_62; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_448 = io_in_dat_mask_63 ? io_in_dat_data_63 : dat_pre_data_63; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_449 = io_in_dat_mask_64 ? io_in_dat_data_64 : dat_pre_data_64; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_450 = io_in_dat_mask_65 ? io_in_dat_data_65 : dat_pre_data_65; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_451 = io_in_dat_mask_66 ? io_in_dat_data_66 : dat_pre_data_66; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_452 = io_in_dat_mask_67 ? io_in_dat_data_67 : dat_pre_data_67; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_453 = io_in_dat_mask_68 ? io_in_dat_data_68 : dat_pre_data_68; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_454 = io_in_dat_mask_69 ? io_in_dat_data_69 : dat_pre_data_69; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_455 = io_in_dat_mask_70 ? io_in_dat_data_70 : dat_pre_data_70; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_456 = io_in_dat_mask_71 ? io_in_dat_data_71 : dat_pre_data_71; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_457 = io_in_dat_mask_72 ? io_in_dat_data_72 : dat_pre_data_72; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_458 = io_in_dat_mask_73 ? io_in_dat_data_73 : dat_pre_data_73; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_459 = io_in_dat_mask_74 ? io_in_dat_data_74 : dat_pre_data_74; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_460 = io_in_dat_mask_75 ? io_in_dat_data_75 : dat_pre_data_75; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_461 = io_in_dat_mask_76 ? io_in_dat_data_76 : dat_pre_data_76; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_462 = io_in_dat_mask_77 ? io_in_dat_data_77 : dat_pre_data_77; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_463 = io_in_dat_mask_78 ? io_in_dat_data_78 : dat_pre_data_78; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_464 = io_in_dat_mask_79 ? io_in_dat_data_79 : dat_pre_data_79; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_465 = io_in_dat_mask_80 ? io_in_dat_data_80 : dat_pre_data_80; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_466 = io_in_dat_mask_81 ? io_in_dat_data_81 : dat_pre_data_81; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_467 = io_in_dat_mask_82 ? io_in_dat_data_82 : dat_pre_data_82; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_468 = io_in_dat_mask_83 ? io_in_dat_data_83 : dat_pre_data_83; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_469 = io_in_dat_mask_84 ? io_in_dat_data_84 : dat_pre_data_84; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_470 = io_in_dat_mask_85 ? io_in_dat_data_85 : dat_pre_data_85; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_471 = io_in_dat_mask_86 ? io_in_dat_data_86 : dat_pre_data_86; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_472 = io_in_dat_mask_87 ? io_in_dat_data_87 : dat_pre_data_87; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_473 = io_in_dat_mask_88 ? io_in_dat_data_88 : dat_pre_data_88; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_474 = io_in_dat_mask_89 ? io_in_dat_data_89 : dat_pre_data_89; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_475 = io_in_dat_mask_90 ? io_in_dat_data_90 : dat_pre_data_90; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_476 = io_in_dat_mask_91 ? io_in_dat_data_91 : dat_pre_data_91; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_477 = io_in_dat_mask_92 ? io_in_dat_data_92 : dat_pre_data_92; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_478 = io_in_dat_mask_93 ? io_in_dat_data_93 : dat_pre_data_93; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_479 = io_in_dat_mask_94 ? io_in_dat_data_94 : dat_pre_data_94; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_480 = io_in_dat_mask_95 ? io_in_dat_data_95 : dat_pre_data_95; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_481 = io_in_dat_mask_96 ? io_in_dat_data_96 : dat_pre_data_96; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_482 = io_in_dat_mask_97 ? io_in_dat_data_97 : dat_pre_data_97; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_483 = io_in_dat_mask_98 ? io_in_dat_data_98 : dat_pre_data_98; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_484 = io_in_dat_mask_99 ? io_in_dat_data_99 : dat_pre_data_99; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_485 = io_in_dat_mask_100 ? io_in_dat_data_100 : dat_pre_data_100; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_486 = io_in_dat_mask_101 ? io_in_dat_data_101 : dat_pre_data_101; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_487 = io_in_dat_mask_102 ? io_in_dat_data_102 : dat_pre_data_102; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_488 = io_in_dat_mask_103 ? io_in_dat_data_103 : dat_pre_data_103; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_489 = io_in_dat_mask_104 ? io_in_dat_data_104 : dat_pre_data_104; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_490 = io_in_dat_mask_105 ? io_in_dat_data_105 : dat_pre_data_105; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_491 = io_in_dat_mask_106 ? io_in_dat_data_106 : dat_pre_data_106; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_492 = io_in_dat_mask_107 ? io_in_dat_data_107 : dat_pre_data_107; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_493 = io_in_dat_mask_108 ? io_in_dat_data_108 : dat_pre_data_108; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_494 = io_in_dat_mask_109 ? io_in_dat_data_109 : dat_pre_data_109; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_495 = io_in_dat_mask_110 ? io_in_dat_data_110 : dat_pre_data_110; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_496 = io_in_dat_mask_111 ? io_in_dat_data_111 : dat_pre_data_111; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_497 = io_in_dat_mask_112 ? io_in_dat_data_112 : dat_pre_data_112; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_498 = io_in_dat_mask_113 ? io_in_dat_data_113 : dat_pre_data_113; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_499 = io_in_dat_mask_114 ? io_in_dat_data_114 : dat_pre_data_114; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_500 = io_in_dat_mask_115 ? io_in_dat_data_115 : dat_pre_data_115; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_501 = io_in_dat_mask_116 ? io_in_dat_data_116 : dat_pre_data_116; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_502 = io_in_dat_mask_117 ? io_in_dat_data_117 : dat_pre_data_117; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_503 = io_in_dat_mask_118 ? io_in_dat_data_118 : dat_pre_data_118; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_504 = io_in_dat_mask_119 ? io_in_dat_data_119 : dat_pre_data_119; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_505 = io_in_dat_mask_120 ? io_in_dat_data_120 : dat_pre_data_120; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_506 = io_in_dat_mask_121 ? io_in_dat_data_121 : dat_pre_data_121; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_507 = io_in_dat_mask_122 ? io_in_dat_data_122 : dat_pre_data_122; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_508 = io_in_dat_mask_123 ? io_in_dat_data_123 : dat_pre_data_123; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_509 = io_in_dat_mask_124 ? io_in_dat_data_124 : dat_pre_data_124; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_510 = io_in_dat_mask_125 ? io_in_dat_data_125 : dat_pre_data_125; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_511 = io_in_dat_mask_126 ? io_in_dat_data_126 : dat_pre_data_126; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_512 = io_in_dat_mask_127 ? io_in_dat_data_127 : dat_pre_data_127; // @[NV_NVDLA_CMAC_CORE_active.scala 92:36]
  assign _GEN_513 = io_in_dat_pvld ? io_in_dat_mask_0 : dat_pre_nz_0; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_514 = io_in_dat_pvld ? io_in_dat_mask_1 : dat_pre_nz_1; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_515 = io_in_dat_pvld ? io_in_dat_mask_2 : dat_pre_nz_2; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_516 = io_in_dat_pvld ? io_in_dat_mask_3 : dat_pre_nz_3; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_517 = io_in_dat_pvld ? io_in_dat_mask_4 : dat_pre_nz_4; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_518 = io_in_dat_pvld ? io_in_dat_mask_5 : dat_pre_nz_5; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_519 = io_in_dat_pvld ? io_in_dat_mask_6 : dat_pre_nz_6; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_520 = io_in_dat_pvld ? io_in_dat_mask_7 : dat_pre_nz_7; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_521 = io_in_dat_pvld ? io_in_dat_mask_8 : dat_pre_nz_8; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_522 = io_in_dat_pvld ? io_in_dat_mask_9 : dat_pre_nz_9; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_523 = io_in_dat_pvld ? io_in_dat_mask_10 : dat_pre_nz_10; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_524 = io_in_dat_pvld ? io_in_dat_mask_11 : dat_pre_nz_11; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_525 = io_in_dat_pvld ? io_in_dat_mask_12 : dat_pre_nz_12; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_526 = io_in_dat_pvld ? io_in_dat_mask_13 : dat_pre_nz_13; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_527 = io_in_dat_pvld ? io_in_dat_mask_14 : dat_pre_nz_14; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_528 = io_in_dat_pvld ? io_in_dat_mask_15 : dat_pre_nz_15; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_529 = io_in_dat_pvld ? io_in_dat_mask_16 : dat_pre_nz_16; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_530 = io_in_dat_pvld ? io_in_dat_mask_17 : dat_pre_nz_17; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_531 = io_in_dat_pvld ? io_in_dat_mask_18 : dat_pre_nz_18; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_532 = io_in_dat_pvld ? io_in_dat_mask_19 : dat_pre_nz_19; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_533 = io_in_dat_pvld ? io_in_dat_mask_20 : dat_pre_nz_20; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_534 = io_in_dat_pvld ? io_in_dat_mask_21 : dat_pre_nz_21; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_535 = io_in_dat_pvld ? io_in_dat_mask_22 : dat_pre_nz_22; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_536 = io_in_dat_pvld ? io_in_dat_mask_23 : dat_pre_nz_23; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_537 = io_in_dat_pvld ? io_in_dat_mask_24 : dat_pre_nz_24; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_538 = io_in_dat_pvld ? io_in_dat_mask_25 : dat_pre_nz_25; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_539 = io_in_dat_pvld ? io_in_dat_mask_26 : dat_pre_nz_26; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_540 = io_in_dat_pvld ? io_in_dat_mask_27 : dat_pre_nz_27; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_541 = io_in_dat_pvld ? io_in_dat_mask_28 : dat_pre_nz_28; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_542 = io_in_dat_pvld ? io_in_dat_mask_29 : dat_pre_nz_29; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_543 = io_in_dat_pvld ? io_in_dat_mask_30 : dat_pre_nz_30; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_544 = io_in_dat_pvld ? io_in_dat_mask_31 : dat_pre_nz_31; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_545 = io_in_dat_pvld ? io_in_dat_mask_32 : dat_pre_nz_32; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_546 = io_in_dat_pvld ? io_in_dat_mask_33 : dat_pre_nz_33; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_547 = io_in_dat_pvld ? io_in_dat_mask_34 : dat_pre_nz_34; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_548 = io_in_dat_pvld ? io_in_dat_mask_35 : dat_pre_nz_35; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_549 = io_in_dat_pvld ? io_in_dat_mask_36 : dat_pre_nz_36; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_550 = io_in_dat_pvld ? io_in_dat_mask_37 : dat_pre_nz_37; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_551 = io_in_dat_pvld ? io_in_dat_mask_38 : dat_pre_nz_38; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_552 = io_in_dat_pvld ? io_in_dat_mask_39 : dat_pre_nz_39; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_553 = io_in_dat_pvld ? io_in_dat_mask_40 : dat_pre_nz_40; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_554 = io_in_dat_pvld ? io_in_dat_mask_41 : dat_pre_nz_41; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_555 = io_in_dat_pvld ? io_in_dat_mask_42 : dat_pre_nz_42; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_556 = io_in_dat_pvld ? io_in_dat_mask_43 : dat_pre_nz_43; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_557 = io_in_dat_pvld ? io_in_dat_mask_44 : dat_pre_nz_44; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_558 = io_in_dat_pvld ? io_in_dat_mask_45 : dat_pre_nz_45; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_559 = io_in_dat_pvld ? io_in_dat_mask_46 : dat_pre_nz_46; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_560 = io_in_dat_pvld ? io_in_dat_mask_47 : dat_pre_nz_47; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_561 = io_in_dat_pvld ? io_in_dat_mask_48 : dat_pre_nz_48; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_562 = io_in_dat_pvld ? io_in_dat_mask_49 : dat_pre_nz_49; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_563 = io_in_dat_pvld ? io_in_dat_mask_50 : dat_pre_nz_50; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_564 = io_in_dat_pvld ? io_in_dat_mask_51 : dat_pre_nz_51; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_565 = io_in_dat_pvld ? io_in_dat_mask_52 : dat_pre_nz_52; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_566 = io_in_dat_pvld ? io_in_dat_mask_53 : dat_pre_nz_53; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_567 = io_in_dat_pvld ? io_in_dat_mask_54 : dat_pre_nz_54; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_568 = io_in_dat_pvld ? io_in_dat_mask_55 : dat_pre_nz_55; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_569 = io_in_dat_pvld ? io_in_dat_mask_56 : dat_pre_nz_56; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_570 = io_in_dat_pvld ? io_in_dat_mask_57 : dat_pre_nz_57; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_571 = io_in_dat_pvld ? io_in_dat_mask_58 : dat_pre_nz_58; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_572 = io_in_dat_pvld ? io_in_dat_mask_59 : dat_pre_nz_59; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_573 = io_in_dat_pvld ? io_in_dat_mask_60 : dat_pre_nz_60; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_574 = io_in_dat_pvld ? io_in_dat_mask_61 : dat_pre_nz_61; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_575 = io_in_dat_pvld ? io_in_dat_mask_62 : dat_pre_nz_62; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_576 = io_in_dat_pvld ? io_in_dat_mask_63 : dat_pre_nz_63; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_577 = io_in_dat_pvld ? io_in_dat_mask_64 : dat_pre_nz_64; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_578 = io_in_dat_pvld ? io_in_dat_mask_65 : dat_pre_nz_65; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_579 = io_in_dat_pvld ? io_in_dat_mask_66 : dat_pre_nz_66; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_580 = io_in_dat_pvld ? io_in_dat_mask_67 : dat_pre_nz_67; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_581 = io_in_dat_pvld ? io_in_dat_mask_68 : dat_pre_nz_68; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_582 = io_in_dat_pvld ? io_in_dat_mask_69 : dat_pre_nz_69; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_583 = io_in_dat_pvld ? io_in_dat_mask_70 : dat_pre_nz_70; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_584 = io_in_dat_pvld ? io_in_dat_mask_71 : dat_pre_nz_71; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_585 = io_in_dat_pvld ? io_in_dat_mask_72 : dat_pre_nz_72; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_586 = io_in_dat_pvld ? io_in_dat_mask_73 : dat_pre_nz_73; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_587 = io_in_dat_pvld ? io_in_dat_mask_74 : dat_pre_nz_74; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_588 = io_in_dat_pvld ? io_in_dat_mask_75 : dat_pre_nz_75; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_589 = io_in_dat_pvld ? io_in_dat_mask_76 : dat_pre_nz_76; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_590 = io_in_dat_pvld ? io_in_dat_mask_77 : dat_pre_nz_77; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_591 = io_in_dat_pvld ? io_in_dat_mask_78 : dat_pre_nz_78; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_592 = io_in_dat_pvld ? io_in_dat_mask_79 : dat_pre_nz_79; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_593 = io_in_dat_pvld ? io_in_dat_mask_80 : dat_pre_nz_80; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_594 = io_in_dat_pvld ? io_in_dat_mask_81 : dat_pre_nz_81; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_595 = io_in_dat_pvld ? io_in_dat_mask_82 : dat_pre_nz_82; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_596 = io_in_dat_pvld ? io_in_dat_mask_83 : dat_pre_nz_83; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_597 = io_in_dat_pvld ? io_in_dat_mask_84 : dat_pre_nz_84; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_598 = io_in_dat_pvld ? io_in_dat_mask_85 : dat_pre_nz_85; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_599 = io_in_dat_pvld ? io_in_dat_mask_86 : dat_pre_nz_86; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_600 = io_in_dat_pvld ? io_in_dat_mask_87 : dat_pre_nz_87; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_601 = io_in_dat_pvld ? io_in_dat_mask_88 : dat_pre_nz_88; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_602 = io_in_dat_pvld ? io_in_dat_mask_89 : dat_pre_nz_89; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_603 = io_in_dat_pvld ? io_in_dat_mask_90 : dat_pre_nz_90; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_604 = io_in_dat_pvld ? io_in_dat_mask_91 : dat_pre_nz_91; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_605 = io_in_dat_pvld ? io_in_dat_mask_92 : dat_pre_nz_92; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_606 = io_in_dat_pvld ? io_in_dat_mask_93 : dat_pre_nz_93; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_607 = io_in_dat_pvld ? io_in_dat_mask_94 : dat_pre_nz_94; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_608 = io_in_dat_pvld ? io_in_dat_mask_95 : dat_pre_nz_95; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_609 = io_in_dat_pvld ? io_in_dat_mask_96 : dat_pre_nz_96; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_610 = io_in_dat_pvld ? io_in_dat_mask_97 : dat_pre_nz_97; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_611 = io_in_dat_pvld ? io_in_dat_mask_98 : dat_pre_nz_98; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_612 = io_in_dat_pvld ? io_in_dat_mask_99 : dat_pre_nz_99; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_613 = io_in_dat_pvld ? io_in_dat_mask_100 : dat_pre_nz_100; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_614 = io_in_dat_pvld ? io_in_dat_mask_101 : dat_pre_nz_101; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_615 = io_in_dat_pvld ? io_in_dat_mask_102 : dat_pre_nz_102; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_616 = io_in_dat_pvld ? io_in_dat_mask_103 : dat_pre_nz_103; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_617 = io_in_dat_pvld ? io_in_dat_mask_104 : dat_pre_nz_104; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_618 = io_in_dat_pvld ? io_in_dat_mask_105 : dat_pre_nz_105; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_619 = io_in_dat_pvld ? io_in_dat_mask_106 : dat_pre_nz_106; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_620 = io_in_dat_pvld ? io_in_dat_mask_107 : dat_pre_nz_107; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_621 = io_in_dat_pvld ? io_in_dat_mask_108 : dat_pre_nz_108; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_622 = io_in_dat_pvld ? io_in_dat_mask_109 : dat_pre_nz_109; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_623 = io_in_dat_pvld ? io_in_dat_mask_110 : dat_pre_nz_110; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_624 = io_in_dat_pvld ? io_in_dat_mask_111 : dat_pre_nz_111; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_625 = io_in_dat_pvld ? io_in_dat_mask_112 : dat_pre_nz_112; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_626 = io_in_dat_pvld ? io_in_dat_mask_113 : dat_pre_nz_113; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_627 = io_in_dat_pvld ? io_in_dat_mask_114 : dat_pre_nz_114; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_628 = io_in_dat_pvld ? io_in_dat_mask_115 : dat_pre_nz_115; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_629 = io_in_dat_pvld ? io_in_dat_mask_116 : dat_pre_nz_116; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_630 = io_in_dat_pvld ? io_in_dat_mask_117 : dat_pre_nz_117; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_631 = io_in_dat_pvld ? io_in_dat_mask_118 : dat_pre_nz_118; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_632 = io_in_dat_pvld ? io_in_dat_mask_119 : dat_pre_nz_119; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_633 = io_in_dat_pvld ? io_in_dat_mask_120 : dat_pre_nz_120; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_634 = io_in_dat_pvld ? io_in_dat_mask_121 : dat_pre_nz_121; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_635 = io_in_dat_pvld ? io_in_dat_mask_122 : dat_pre_nz_122; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_636 = io_in_dat_pvld ? io_in_dat_mask_123 : dat_pre_nz_123; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_637 = io_in_dat_pvld ? io_in_dat_mask_124 : dat_pre_nz_124; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_638 = io_in_dat_pvld ? io_in_dat_mask_125 : dat_pre_nz_125; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_639 = io_in_dat_pvld ? io_in_dat_mask_126 : dat_pre_nz_126; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_640 = io_in_dat_pvld ? io_in_dat_mask_127 : dat_pre_nz_127; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_769 = io_in_dat_pvld ? io_in_dat_stripe_st : dat_pre_stripe_st_out_0; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _GEN_770 = io_in_dat_pvld ? io_in_dat_stripe_end : dat_pre_stripe_end_out_0; // @[NV_NVDLA_CMAC_CORE_active.scala 89:25]
  assign _T_27793 = dat_pre_stripe_st_out_0 ? 1'h0 : wt_sd_pvld_0; // @[NV_NVDLA_CMAC_CORE_active.scala 115:58]
  assign wt_sd_pvld_w_0 = wt_pre_sel_0 ? 1'h1 : _T_27793; // @[NV_NVDLA_CMAC_CORE_active.scala 115:31]
  assign _GEN_771 = wt_pre_nz_0 ? wt_pre_data_0 : wt_sd_data_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_772 = wt_pre_nz_1 ? wt_pre_data_1 : wt_sd_data_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_773 = wt_pre_nz_2 ? wt_pre_data_2 : wt_sd_data_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_774 = wt_pre_nz_3 ? wt_pre_data_3 : wt_sd_data_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_775 = wt_pre_nz_4 ? wt_pre_data_4 : wt_sd_data_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_776 = wt_pre_nz_5 ? wt_pre_data_5 : wt_sd_data_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_777 = wt_pre_nz_6 ? wt_pre_data_6 : wt_sd_data_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_778 = wt_pre_nz_7 ? wt_pre_data_7 : wt_sd_data_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_779 = wt_pre_nz_8 ? wt_pre_data_8 : wt_sd_data_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_780 = wt_pre_nz_9 ? wt_pre_data_9 : wt_sd_data_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_781 = wt_pre_nz_10 ? wt_pre_data_10 : wt_sd_data_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_782 = wt_pre_nz_11 ? wt_pre_data_11 : wt_sd_data_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_783 = wt_pre_nz_12 ? wt_pre_data_12 : wt_sd_data_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_784 = wt_pre_nz_13 ? wt_pre_data_13 : wt_sd_data_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_785 = wt_pre_nz_14 ? wt_pre_data_14 : wt_sd_data_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_786 = wt_pre_nz_15 ? wt_pre_data_15 : wt_sd_data_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_787 = wt_pre_nz_16 ? wt_pre_data_16 : wt_sd_data_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_788 = wt_pre_nz_17 ? wt_pre_data_17 : wt_sd_data_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_789 = wt_pre_nz_18 ? wt_pre_data_18 : wt_sd_data_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_790 = wt_pre_nz_19 ? wt_pre_data_19 : wt_sd_data_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_791 = wt_pre_nz_20 ? wt_pre_data_20 : wt_sd_data_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_792 = wt_pre_nz_21 ? wt_pre_data_21 : wt_sd_data_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_793 = wt_pre_nz_22 ? wt_pre_data_22 : wt_sd_data_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_794 = wt_pre_nz_23 ? wt_pre_data_23 : wt_sd_data_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_795 = wt_pre_nz_24 ? wt_pre_data_24 : wt_sd_data_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_796 = wt_pre_nz_25 ? wt_pre_data_25 : wt_sd_data_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_797 = wt_pre_nz_26 ? wt_pre_data_26 : wt_sd_data_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_798 = wt_pre_nz_27 ? wt_pre_data_27 : wt_sd_data_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_799 = wt_pre_nz_28 ? wt_pre_data_28 : wt_sd_data_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_800 = wt_pre_nz_29 ? wt_pre_data_29 : wt_sd_data_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_801 = wt_pre_nz_30 ? wt_pre_data_30 : wt_sd_data_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_802 = wt_pre_nz_31 ? wt_pre_data_31 : wt_sd_data_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_803 = wt_pre_nz_32 ? wt_pre_data_32 : wt_sd_data_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_804 = wt_pre_nz_33 ? wt_pre_data_33 : wt_sd_data_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_805 = wt_pre_nz_34 ? wt_pre_data_34 : wt_sd_data_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_806 = wt_pre_nz_35 ? wt_pre_data_35 : wt_sd_data_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_807 = wt_pre_nz_36 ? wt_pre_data_36 : wt_sd_data_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_808 = wt_pre_nz_37 ? wt_pre_data_37 : wt_sd_data_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_809 = wt_pre_nz_38 ? wt_pre_data_38 : wt_sd_data_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_810 = wt_pre_nz_39 ? wt_pre_data_39 : wt_sd_data_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_811 = wt_pre_nz_40 ? wt_pre_data_40 : wt_sd_data_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_812 = wt_pre_nz_41 ? wt_pre_data_41 : wt_sd_data_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_813 = wt_pre_nz_42 ? wt_pre_data_42 : wt_sd_data_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_814 = wt_pre_nz_43 ? wt_pre_data_43 : wt_sd_data_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_815 = wt_pre_nz_44 ? wt_pre_data_44 : wt_sd_data_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_816 = wt_pre_nz_45 ? wt_pre_data_45 : wt_sd_data_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_817 = wt_pre_nz_46 ? wt_pre_data_46 : wt_sd_data_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_818 = wt_pre_nz_47 ? wt_pre_data_47 : wt_sd_data_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_819 = wt_pre_nz_48 ? wt_pre_data_48 : wt_sd_data_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_820 = wt_pre_nz_49 ? wt_pre_data_49 : wt_sd_data_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_821 = wt_pre_nz_50 ? wt_pre_data_50 : wt_sd_data_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_822 = wt_pre_nz_51 ? wt_pre_data_51 : wt_sd_data_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_823 = wt_pre_nz_52 ? wt_pre_data_52 : wt_sd_data_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_824 = wt_pre_nz_53 ? wt_pre_data_53 : wt_sd_data_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_825 = wt_pre_nz_54 ? wt_pre_data_54 : wt_sd_data_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_826 = wt_pre_nz_55 ? wt_pre_data_55 : wt_sd_data_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_827 = wt_pre_nz_56 ? wt_pre_data_56 : wt_sd_data_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_828 = wt_pre_nz_57 ? wt_pre_data_57 : wt_sd_data_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_829 = wt_pre_nz_58 ? wt_pre_data_58 : wt_sd_data_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_830 = wt_pre_nz_59 ? wt_pre_data_59 : wt_sd_data_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_831 = wt_pre_nz_60 ? wt_pre_data_60 : wt_sd_data_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_832 = wt_pre_nz_61 ? wt_pre_data_61 : wt_sd_data_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_833 = wt_pre_nz_62 ? wt_pre_data_62 : wt_sd_data_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_834 = wt_pre_nz_63 ? wt_pre_data_63 : wt_sd_data_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_835 = wt_pre_nz_64 ? wt_pre_data_64 : wt_sd_data_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_836 = wt_pre_nz_65 ? wt_pre_data_65 : wt_sd_data_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_837 = wt_pre_nz_66 ? wt_pre_data_66 : wt_sd_data_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_838 = wt_pre_nz_67 ? wt_pre_data_67 : wt_sd_data_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_839 = wt_pre_nz_68 ? wt_pre_data_68 : wt_sd_data_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_840 = wt_pre_nz_69 ? wt_pre_data_69 : wt_sd_data_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_841 = wt_pre_nz_70 ? wt_pre_data_70 : wt_sd_data_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_842 = wt_pre_nz_71 ? wt_pre_data_71 : wt_sd_data_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_843 = wt_pre_nz_72 ? wt_pre_data_72 : wt_sd_data_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_844 = wt_pre_nz_73 ? wt_pre_data_73 : wt_sd_data_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_845 = wt_pre_nz_74 ? wt_pre_data_74 : wt_sd_data_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_846 = wt_pre_nz_75 ? wt_pre_data_75 : wt_sd_data_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_847 = wt_pre_nz_76 ? wt_pre_data_76 : wt_sd_data_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_848 = wt_pre_nz_77 ? wt_pre_data_77 : wt_sd_data_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_849 = wt_pre_nz_78 ? wt_pre_data_78 : wt_sd_data_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_850 = wt_pre_nz_79 ? wt_pre_data_79 : wt_sd_data_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_851 = wt_pre_nz_80 ? wt_pre_data_80 : wt_sd_data_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_852 = wt_pre_nz_81 ? wt_pre_data_81 : wt_sd_data_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_853 = wt_pre_nz_82 ? wt_pre_data_82 : wt_sd_data_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_854 = wt_pre_nz_83 ? wt_pre_data_83 : wt_sd_data_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_855 = wt_pre_nz_84 ? wt_pre_data_84 : wt_sd_data_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_856 = wt_pre_nz_85 ? wt_pre_data_85 : wt_sd_data_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_857 = wt_pre_nz_86 ? wt_pre_data_86 : wt_sd_data_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_858 = wt_pre_nz_87 ? wt_pre_data_87 : wt_sd_data_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_859 = wt_pre_nz_88 ? wt_pre_data_88 : wt_sd_data_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_860 = wt_pre_nz_89 ? wt_pre_data_89 : wt_sd_data_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_861 = wt_pre_nz_90 ? wt_pre_data_90 : wt_sd_data_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_862 = wt_pre_nz_91 ? wt_pre_data_91 : wt_sd_data_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_863 = wt_pre_nz_92 ? wt_pre_data_92 : wt_sd_data_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_864 = wt_pre_nz_93 ? wt_pre_data_93 : wt_sd_data_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_865 = wt_pre_nz_94 ? wt_pre_data_94 : wt_sd_data_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_866 = wt_pre_nz_95 ? wt_pre_data_95 : wt_sd_data_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_867 = wt_pre_nz_96 ? wt_pre_data_96 : wt_sd_data_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_868 = wt_pre_nz_97 ? wt_pre_data_97 : wt_sd_data_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_869 = wt_pre_nz_98 ? wt_pre_data_98 : wt_sd_data_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_870 = wt_pre_nz_99 ? wt_pre_data_99 : wt_sd_data_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_871 = wt_pre_nz_100 ? wt_pre_data_100 : wt_sd_data_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_872 = wt_pre_nz_101 ? wt_pre_data_101 : wt_sd_data_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_873 = wt_pre_nz_102 ? wt_pre_data_102 : wt_sd_data_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_874 = wt_pre_nz_103 ? wt_pre_data_103 : wt_sd_data_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_875 = wt_pre_nz_104 ? wt_pre_data_104 : wt_sd_data_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_876 = wt_pre_nz_105 ? wt_pre_data_105 : wt_sd_data_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_877 = wt_pre_nz_106 ? wt_pre_data_106 : wt_sd_data_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_878 = wt_pre_nz_107 ? wt_pre_data_107 : wt_sd_data_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_879 = wt_pre_nz_108 ? wt_pre_data_108 : wt_sd_data_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_880 = wt_pre_nz_109 ? wt_pre_data_109 : wt_sd_data_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_881 = wt_pre_nz_110 ? wt_pre_data_110 : wt_sd_data_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_882 = wt_pre_nz_111 ? wt_pre_data_111 : wt_sd_data_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_883 = wt_pre_nz_112 ? wt_pre_data_112 : wt_sd_data_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_884 = wt_pre_nz_113 ? wt_pre_data_113 : wt_sd_data_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_885 = wt_pre_nz_114 ? wt_pre_data_114 : wt_sd_data_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_886 = wt_pre_nz_115 ? wt_pre_data_115 : wt_sd_data_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_887 = wt_pre_nz_116 ? wt_pre_data_116 : wt_sd_data_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_888 = wt_pre_nz_117 ? wt_pre_data_117 : wt_sd_data_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_889 = wt_pre_nz_118 ? wt_pre_data_118 : wt_sd_data_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_890 = wt_pre_nz_119 ? wt_pre_data_119 : wt_sd_data_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_891 = wt_pre_nz_120 ? wt_pre_data_120 : wt_sd_data_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_892 = wt_pre_nz_121 ? wt_pre_data_121 : wt_sd_data_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_893 = wt_pre_nz_122 ? wt_pre_data_122 : wt_sd_data_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_894 = wt_pre_nz_123 ? wt_pre_data_123 : wt_sd_data_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_895 = wt_pre_nz_124 ? wt_pre_data_124 : wt_sd_data_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_896 = wt_pre_nz_125 ? wt_pre_data_125 : wt_sd_data_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_897 = wt_pre_nz_126 ? wt_pre_data_126 : wt_sd_data_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_898 = wt_pre_nz_127 ? wt_pre_data_127 : wt_sd_data_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 120:35]
  assign _GEN_899 = wt_pre_sel_0 ? wt_pre_nz_0 : wt_sd_nz_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_900 = wt_pre_sel_0 ? wt_pre_nz_1 : wt_sd_nz_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_901 = wt_pre_sel_0 ? wt_pre_nz_2 : wt_sd_nz_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_902 = wt_pre_sel_0 ? wt_pre_nz_3 : wt_sd_nz_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_903 = wt_pre_sel_0 ? wt_pre_nz_4 : wt_sd_nz_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_904 = wt_pre_sel_0 ? wt_pre_nz_5 : wt_sd_nz_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_905 = wt_pre_sel_0 ? wt_pre_nz_6 : wt_sd_nz_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_906 = wt_pre_sel_0 ? wt_pre_nz_7 : wt_sd_nz_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_907 = wt_pre_sel_0 ? wt_pre_nz_8 : wt_sd_nz_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_908 = wt_pre_sel_0 ? wt_pre_nz_9 : wt_sd_nz_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_909 = wt_pre_sel_0 ? wt_pre_nz_10 : wt_sd_nz_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_910 = wt_pre_sel_0 ? wt_pre_nz_11 : wt_sd_nz_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_911 = wt_pre_sel_0 ? wt_pre_nz_12 : wt_sd_nz_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_912 = wt_pre_sel_0 ? wt_pre_nz_13 : wt_sd_nz_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_913 = wt_pre_sel_0 ? wt_pre_nz_14 : wt_sd_nz_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_914 = wt_pre_sel_0 ? wt_pre_nz_15 : wt_sd_nz_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_915 = wt_pre_sel_0 ? wt_pre_nz_16 : wt_sd_nz_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_916 = wt_pre_sel_0 ? wt_pre_nz_17 : wt_sd_nz_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_917 = wt_pre_sel_0 ? wt_pre_nz_18 : wt_sd_nz_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_918 = wt_pre_sel_0 ? wt_pre_nz_19 : wt_sd_nz_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_919 = wt_pre_sel_0 ? wt_pre_nz_20 : wt_sd_nz_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_920 = wt_pre_sel_0 ? wt_pre_nz_21 : wt_sd_nz_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_921 = wt_pre_sel_0 ? wt_pre_nz_22 : wt_sd_nz_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_922 = wt_pre_sel_0 ? wt_pre_nz_23 : wt_sd_nz_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_923 = wt_pre_sel_0 ? wt_pre_nz_24 : wt_sd_nz_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_924 = wt_pre_sel_0 ? wt_pre_nz_25 : wt_sd_nz_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_925 = wt_pre_sel_0 ? wt_pre_nz_26 : wt_sd_nz_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_926 = wt_pre_sel_0 ? wt_pre_nz_27 : wt_sd_nz_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_927 = wt_pre_sel_0 ? wt_pre_nz_28 : wt_sd_nz_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_928 = wt_pre_sel_0 ? wt_pre_nz_29 : wt_sd_nz_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_929 = wt_pre_sel_0 ? wt_pre_nz_30 : wt_sd_nz_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_930 = wt_pre_sel_0 ? wt_pre_nz_31 : wt_sd_nz_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_931 = wt_pre_sel_0 ? wt_pre_nz_32 : wt_sd_nz_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_932 = wt_pre_sel_0 ? wt_pre_nz_33 : wt_sd_nz_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_933 = wt_pre_sel_0 ? wt_pre_nz_34 : wt_sd_nz_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_934 = wt_pre_sel_0 ? wt_pre_nz_35 : wt_sd_nz_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_935 = wt_pre_sel_0 ? wt_pre_nz_36 : wt_sd_nz_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_936 = wt_pre_sel_0 ? wt_pre_nz_37 : wt_sd_nz_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_937 = wt_pre_sel_0 ? wt_pre_nz_38 : wt_sd_nz_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_938 = wt_pre_sel_0 ? wt_pre_nz_39 : wt_sd_nz_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_939 = wt_pre_sel_0 ? wt_pre_nz_40 : wt_sd_nz_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_940 = wt_pre_sel_0 ? wt_pre_nz_41 : wt_sd_nz_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_941 = wt_pre_sel_0 ? wt_pre_nz_42 : wt_sd_nz_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_942 = wt_pre_sel_0 ? wt_pre_nz_43 : wt_sd_nz_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_943 = wt_pre_sel_0 ? wt_pre_nz_44 : wt_sd_nz_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_944 = wt_pre_sel_0 ? wt_pre_nz_45 : wt_sd_nz_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_945 = wt_pre_sel_0 ? wt_pre_nz_46 : wt_sd_nz_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_946 = wt_pre_sel_0 ? wt_pre_nz_47 : wt_sd_nz_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_947 = wt_pre_sel_0 ? wt_pre_nz_48 : wt_sd_nz_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_948 = wt_pre_sel_0 ? wt_pre_nz_49 : wt_sd_nz_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_949 = wt_pre_sel_0 ? wt_pre_nz_50 : wt_sd_nz_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_950 = wt_pre_sel_0 ? wt_pre_nz_51 : wt_sd_nz_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_951 = wt_pre_sel_0 ? wt_pre_nz_52 : wt_sd_nz_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_952 = wt_pre_sel_0 ? wt_pre_nz_53 : wt_sd_nz_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_953 = wt_pre_sel_0 ? wt_pre_nz_54 : wt_sd_nz_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_954 = wt_pre_sel_0 ? wt_pre_nz_55 : wt_sd_nz_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_955 = wt_pre_sel_0 ? wt_pre_nz_56 : wt_sd_nz_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_956 = wt_pre_sel_0 ? wt_pre_nz_57 : wt_sd_nz_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_957 = wt_pre_sel_0 ? wt_pre_nz_58 : wt_sd_nz_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_958 = wt_pre_sel_0 ? wt_pre_nz_59 : wt_sd_nz_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_959 = wt_pre_sel_0 ? wt_pre_nz_60 : wt_sd_nz_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_960 = wt_pre_sel_0 ? wt_pre_nz_61 : wt_sd_nz_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_961 = wt_pre_sel_0 ? wt_pre_nz_62 : wt_sd_nz_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_962 = wt_pre_sel_0 ? wt_pre_nz_63 : wt_sd_nz_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_963 = wt_pre_sel_0 ? wt_pre_nz_64 : wt_sd_nz_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_964 = wt_pre_sel_0 ? wt_pre_nz_65 : wt_sd_nz_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_965 = wt_pre_sel_0 ? wt_pre_nz_66 : wt_sd_nz_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_966 = wt_pre_sel_0 ? wt_pre_nz_67 : wt_sd_nz_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_967 = wt_pre_sel_0 ? wt_pre_nz_68 : wt_sd_nz_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_968 = wt_pre_sel_0 ? wt_pre_nz_69 : wt_sd_nz_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_969 = wt_pre_sel_0 ? wt_pre_nz_70 : wt_sd_nz_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_970 = wt_pre_sel_0 ? wt_pre_nz_71 : wt_sd_nz_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_971 = wt_pre_sel_0 ? wt_pre_nz_72 : wt_sd_nz_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_972 = wt_pre_sel_0 ? wt_pre_nz_73 : wt_sd_nz_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_973 = wt_pre_sel_0 ? wt_pre_nz_74 : wt_sd_nz_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_974 = wt_pre_sel_0 ? wt_pre_nz_75 : wt_sd_nz_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_975 = wt_pre_sel_0 ? wt_pre_nz_76 : wt_sd_nz_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_976 = wt_pre_sel_0 ? wt_pre_nz_77 : wt_sd_nz_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_977 = wt_pre_sel_0 ? wt_pre_nz_78 : wt_sd_nz_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_978 = wt_pre_sel_0 ? wt_pre_nz_79 : wt_sd_nz_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_979 = wt_pre_sel_0 ? wt_pre_nz_80 : wt_sd_nz_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_980 = wt_pre_sel_0 ? wt_pre_nz_81 : wt_sd_nz_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_981 = wt_pre_sel_0 ? wt_pre_nz_82 : wt_sd_nz_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_982 = wt_pre_sel_0 ? wt_pre_nz_83 : wt_sd_nz_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_983 = wt_pre_sel_0 ? wt_pre_nz_84 : wt_sd_nz_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_984 = wt_pre_sel_0 ? wt_pre_nz_85 : wt_sd_nz_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_985 = wt_pre_sel_0 ? wt_pre_nz_86 : wt_sd_nz_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_986 = wt_pre_sel_0 ? wt_pre_nz_87 : wt_sd_nz_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_987 = wt_pre_sel_0 ? wt_pre_nz_88 : wt_sd_nz_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_988 = wt_pre_sel_0 ? wt_pre_nz_89 : wt_sd_nz_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_989 = wt_pre_sel_0 ? wt_pre_nz_90 : wt_sd_nz_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_990 = wt_pre_sel_0 ? wt_pre_nz_91 : wt_sd_nz_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_991 = wt_pre_sel_0 ? wt_pre_nz_92 : wt_sd_nz_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_992 = wt_pre_sel_0 ? wt_pre_nz_93 : wt_sd_nz_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_993 = wt_pre_sel_0 ? wt_pre_nz_94 : wt_sd_nz_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_994 = wt_pre_sel_0 ? wt_pre_nz_95 : wt_sd_nz_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_995 = wt_pre_sel_0 ? wt_pre_nz_96 : wt_sd_nz_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_996 = wt_pre_sel_0 ? wt_pre_nz_97 : wt_sd_nz_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_997 = wt_pre_sel_0 ? wt_pre_nz_98 : wt_sd_nz_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_998 = wt_pre_sel_0 ? wt_pre_nz_99 : wt_sd_nz_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_999 = wt_pre_sel_0 ? wt_pre_nz_100 : wt_sd_nz_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1000 = wt_pre_sel_0 ? wt_pre_nz_101 : wt_sd_nz_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1001 = wt_pre_sel_0 ? wt_pre_nz_102 : wt_sd_nz_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1002 = wt_pre_sel_0 ? wt_pre_nz_103 : wt_sd_nz_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1003 = wt_pre_sel_0 ? wt_pre_nz_104 : wt_sd_nz_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1004 = wt_pre_sel_0 ? wt_pre_nz_105 : wt_sd_nz_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1005 = wt_pre_sel_0 ? wt_pre_nz_106 : wt_sd_nz_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1006 = wt_pre_sel_0 ? wt_pre_nz_107 : wt_sd_nz_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1007 = wt_pre_sel_0 ? wt_pre_nz_108 : wt_sd_nz_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1008 = wt_pre_sel_0 ? wt_pre_nz_109 : wt_sd_nz_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1009 = wt_pre_sel_0 ? wt_pre_nz_110 : wt_sd_nz_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1010 = wt_pre_sel_0 ? wt_pre_nz_111 : wt_sd_nz_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1011 = wt_pre_sel_0 ? wt_pre_nz_112 : wt_sd_nz_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1012 = wt_pre_sel_0 ? wt_pre_nz_113 : wt_sd_nz_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1013 = wt_pre_sel_0 ? wt_pre_nz_114 : wt_sd_nz_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1014 = wt_pre_sel_0 ? wt_pre_nz_115 : wt_sd_nz_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1015 = wt_pre_sel_0 ? wt_pre_nz_116 : wt_sd_nz_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1016 = wt_pre_sel_0 ? wt_pre_nz_117 : wt_sd_nz_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1017 = wt_pre_sel_0 ? wt_pre_nz_118 : wt_sd_nz_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1018 = wt_pre_sel_0 ? wt_pre_nz_119 : wt_sd_nz_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1019 = wt_pre_sel_0 ? wt_pre_nz_120 : wt_sd_nz_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1020 = wt_pre_sel_0 ? wt_pre_nz_121 : wt_sd_nz_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1021 = wt_pre_sel_0 ? wt_pre_nz_122 : wt_sd_nz_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1022 = wt_pre_sel_0 ? wt_pre_nz_123 : wt_sd_nz_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1023 = wt_pre_sel_0 ? wt_pre_nz_124 : wt_sd_nz_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1024 = wt_pre_sel_0 ? wt_pre_nz_125 : wt_sd_nz_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1025 = wt_pre_sel_0 ? wt_pre_nz_126 : wt_sd_nz_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _GEN_1026 = wt_pre_sel_0 ? wt_pre_nz_127 : wt_sd_nz_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 117:28]
  assign _T_50631 = dat_actv_stripe_end_0 ? 1'h0 : wt_actv_vld_0; // @[NV_NVDLA_CMAC_CORE_active.scala 141:78]
  assign wt_actv_pvld_w_0 = dat_pre_stripe_st_out_0 ? wt_sd_pvld_0 : _T_50631; // @[NV_NVDLA_CMAC_CORE_active.scala 141:33]
  assign _T_50633 = dat_pre_stripe_st_out_0 & wt_actv_pvld_w_0; // @[NV_NVDLA_CMAC_CORE_active.scala 145:42]
  assign _GEN_1155 = wt_sd_nz_0_0 ? wt_sd_data_0_0 : wt_actv_data_out_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1156 = _T_50633 ? wt_sd_nz_0_0 : wt_actv_nz_out_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1158 = wt_sd_nz_0_1 ? wt_sd_data_0_1 : wt_actv_data_out_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1159 = _T_50633 ? wt_sd_nz_0_1 : wt_actv_nz_out_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1161 = wt_sd_nz_0_2 ? wt_sd_data_0_2 : wt_actv_data_out_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1162 = _T_50633 ? wt_sd_nz_0_2 : wt_actv_nz_out_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1164 = wt_sd_nz_0_3 ? wt_sd_data_0_3 : wt_actv_data_out_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1165 = _T_50633 ? wt_sd_nz_0_3 : wt_actv_nz_out_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1167 = wt_sd_nz_0_4 ? wt_sd_data_0_4 : wt_actv_data_out_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1168 = _T_50633 ? wt_sd_nz_0_4 : wt_actv_nz_out_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1170 = wt_sd_nz_0_5 ? wt_sd_data_0_5 : wt_actv_data_out_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1171 = _T_50633 ? wt_sd_nz_0_5 : wt_actv_nz_out_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1173 = wt_sd_nz_0_6 ? wt_sd_data_0_6 : wt_actv_data_out_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1174 = _T_50633 ? wt_sd_nz_0_6 : wt_actv_nz_out_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1176 = wt_sd_nz_0_7 ? wt_sd_data_0_7 : wt_actv_data_out_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1177 = _T_50633 ? wt_sd_nz_0_7 : wt_actv_nz_out_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1179 = wt_sd_nz_0_8 ? wt_sd_data_0_8 : wt_actv_data_out_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1180 = _T_50633 ? wt_sd_nz_0_8 : wt_actv_nz_out_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1182 = wt_sd_nz_0_9 ? wt_sd_data_0_9 : wt_actv_data_out_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1183 = _T_50633 ? wt_sd_nz_0_9 : wt_actv_nz_out_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1185 = wt_sd_nz_0_10 ? wt_sd_data_0_10 : wt_actv_data_out_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1186 = _T_50633 ? wt_sd_nz_0_10 : wt_actv_nz_out_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1188 = wt_sd_nz_0_11 ? wt_sd_data_0_11 : wt_actv_data_out_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1189 = _T_50633 ? wt_sd_nz_0_11 : wt_actv_nz_out_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1191 = wt_sd_nz_0_12 ? wt_sd_data_0_12 : wt_actv_data_out_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1192 = _T_50633 ? wt_sd_nz_0_12 : wt_actv_nz_out_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1194 = wt_sd_nz_0_13 ? wt_sd_data_0_13 : wt_actv_data_out_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1195 = _T_50633 ? wt_sd_nz_0_13 : wt_actv_nz_out_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1197 = wt_sd_nz_0_14 ? wt_sd_data_0_14 : wt_actv_data_out_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1198 = _T_50633 ? wt_sd_nz_0_14 : wt_actv_nz_out_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1200 = wt_sd_nz_0_15 ? wt_sd_data_0_15 : wt_actv_data_out_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1201 = _T_50633 ? wt_sd_nz_0_15 : wt_actv_nz_out_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1203 = wt_sd_nz_0_16 ? wt_sd_data_0_16 : wt_actv_data_out_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1204 = _T_50633 ? wt_sd_nz_0_16 : wt_actv_nz_out_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1206 = wt_sd_nz_0_17 ? wt_sd_data_0_17 : wt_actv_data_out_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1207 = _T_50633 ? wt_sd_nz_0_17 : wt_actv_nz_out_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1209 = wt_sd_nz_0_18 ? wt_sd_data_0_18 : wt_actv_data_out_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1210 = _T_50633 ? wt_sd_nz_0_18 : wt_actv_nz_out_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1212 = wt_sd_nz_0_19 ? wt_sd_data_0_19 : wt_actv_data_out_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1213 = _T_50633 ? wt_sd_nz_0_19 : wt_actv_nz_out_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1215 = wt_sd_nz_0_20 ? wt_sd_data_0_20 : wt_actv_data_out_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1216 = _T_50633 ? wt_sd_nz_0_20 : wt_actv_nz_out_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1218 = wt_sd_nz_0_21 ? wt_sd_data_0_21 : wt_actv_data_out_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1219 = _T_50633 ? wt_sd_nz_0_21 : wt_actv_nz_out_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1221 = wt_sd_nz_0_22 ? wt_sd_data_0_22 : wt_actv_data_out_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1222 = _T_50633 ? wt_sd_nz_0_22 : wt_actv_nz_out_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1224 = wt_sd_nz_0_23 ? wt_sd_data_0_23 : wt_actv_data_out_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1225 = _T_50633 ? wt_sd_nz_0_23 : wt_actv_nz_out_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1227 = wt_sd_nz_0_24 ? wt_sd_data_0_24 : wt_actv_data_out_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1228 = _T_50633 ? wt_sd_nz_0_24 : wt_actv_nz_out_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1230 = wt_sd_nz_0_25 ? wt_sd_data_0_25 : wt_actv_data_out_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1231 = _T_50633 ? wt_sd_nz_0_25 : wt_actv_nz_out_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1233 = wt_sd_nz_0_26 ? wt_sd_data_0_26 : wt_actv_data_out_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1234 = _T_50633 ? wt_sd_nz_0_26 : wt_actv_nz_out_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1236 = wt_sd_nz_0_27 ? wt_sd_data_0_27 : wt_actv_data_out_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1237 = _T_50633 ? wt_sd_nz_0_27 : wt_actv_nz_out_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1239 = wt_sd_nz_0_28 ? wt_sd_data_0_28 : wt_actv_data_out_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1240 = _T_50633 ? wt_sd_nz_0_28 : wt_actv_nz_out_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1242 = wt_sd_nz_0_29 ? wt_sd_data_0_29 : wt_actv_data_out_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1243 = _T_50633 ? wt_sd_nz_0_29 : wt_actv_nz_out_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1245 = wt_sd_nz_0_30 ? wt_sd_data_0_30 : wt_actv_data_out_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1246 = _T_50633 ? wt_sd_nz_0_30 : wt_actv_nz_out_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1248 = wt_sd_nz_0_31 ? wt_sd_data_0_31 : wt_actv_data_out_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1249 = _T_50633 ? wt_sd_nz_0_31 : wt_actv_nz_out_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1251 = wt_sd_nz_0_32 ? wt_sd_data_0_32 : wt_actv_data_out_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1252 = _T_50633 ? wt_sd_nz_0_32 : wt_actv_nz_out_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1254 = wt_sd_nz_0_33 ? wt_sd_data_0_33 : wt_actv_data_out_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1255 = _T_50633 ? wt_sd_nz_0_33 : wt_actv_nz_out_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1257 = wt_sd_nz_0_34 ? wt_sd_data_0_34 : wt_actv_data_out_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1258 = _T_50633 ? wt_sd_nz_0_34 : wt_actv_nz_out_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1260 = wt_sd_nz_0_35 ? wt_sd_data_0_35 : wt_actv_data_out_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1261 = _T_50633 ? wt_sd_nz_0_35 : wt_actv_nz_out_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1263 = wt_sd_nz_0_36 ? wt_sd_data_0_36 : wt_actv_data_out_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1264 = _T_50633 ? wt_sd_nz_0_36 : wt_actv_nz_out_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1266 = wt_sd_nz_0_37 ? wt_sd_data_0_37 : wt_actv_data_out_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1267 = _T_50633 ? wt_sd_nz_0_37 : wt_actv_nz_out_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1269 = wt_sd_nz_0_38 ? wt_sd_data_0_38 : wt_actv_data_out_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1270 = _T_50633 ? wt_sd_nz_0_38 : wt_actv_nz_out_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1272 = wt_sd_nz_0_39 ? wt_sd_data_0_39 : wt_actv_data_out_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1273 = _T_50633 ? wt_sd_nz_0_39 : wt_actv_nz_out_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1275 = wt_sd_nz_0_40 ? wt_sd_data_0_40 : wt_actv_data_out_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1276 = _T_50633 ? wt_sd_nz_0_40 : wt_actv_nz_out_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1278 = wt_sd_nz_0_41 ? wt_sd_data_0_41 : wt_actv_data_out_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1279 = _T_50633 ? wt_sd_nz_0_41 : wt_actv_nz_out_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1281 = wt_sd_nz_0_42 ? wt_sd_data_0_42 : wt_actv_data_out_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1282 = _T_50633 ? wt_sd_nz_0_42 : wt_actv_nz_out_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1284 = wt_sd_nz_0_43 ? wt_sd_data_0_43 : wt_actv_data_out_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1285 = _T_50633 ? wt_sd_nz_0_43 : wt_actv_nz_out_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1287 = wt_sd_nz_0_44 ? wt_sd_data_0_44 : wt_actv_data_out_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1288 = _T_50633 ? wt_sd_nz_0_44 : wt_actv_nz_out_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1290 = wt_sd_nz_0_45 ? wt_sd_data_0_45 : wt_actv_data_out_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1291 = _T_50633 ? wt_sd_nz_0_45 : wt_actv_nz_out_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1293 = wt_sd_nz_0_46 ? wt_sd_data_0_46 : wt_actv_data_out_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1294 = _T_50633 ? wt_sd_nz_0_46 : wt_actv_nz_out_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1296 = wt_sd_nz_0_47 ? wt_sd_data_0_47 : wt_actv_data_out_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1297 = _T_50633 ? wt_sd_nz_0_47 : wt_actv_nz_out_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1299 = wt_sd_nz_0_48 ? wt_sd_data_0_48 : wt_actv_data_out_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1300 = _T_50633 ? wt_sd_nz_0_48 : wt_actv_nz_out_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1302 = wt_sd_nz_0_49 ? wt_sd_data_0_49 : wt_actv_data_out_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1303 = _T_50633 ? wt_sd_nz_0_49 : wt_actv_nz_out_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1305 = wt_sd_nz_0_50 ? wt_sd_data_0_50 : wt_actv_data_out_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1306 = _T_50633 ? wt_sd_nz_0_50 : wt_actv_nz_out_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1308 = wt_sd_nz_0_51 ? wt_sd_data_0_51 : wt_actv_data_out_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1309 = _T_50633 ? wt_sd_nz_0_51 : wt_actv_nz_out_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1311 = wt_sd_nz_0_52 ? wt_sd_data_0_52 : wt_actv_data_out_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1312 = _T_50633 ? wt_sd_nz_0_52 : wt_actv_nz_out_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1314 = wt_sd_nz_0_53 ? wt_sd_data_0_53 : wt_actv_data_out_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1315 = _T_50633 ? wt_sd_nz_0_53 : wt_actv_nz_out_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1317 = wt_sd_nz_0_54 ? wt_sd_data_0_54 : wt_actv_data_out_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1318 = _T_50633 ? wt_sd_nz_0_54 : wt_actv_nz_out_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1320 = wt_sd_nz_0_55 ? wt_sd_data_0_55 : wt_actv_data_out_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1321 = _T_50633 ? wt_sd_nz_0_55 : wt_actv_nz_out_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1323 = wt_sd_nz_0_56 ? wt_sd_data_0_56 : wt_actv_data_out_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1324 = _T_50633 ? wt_sd_nz_0_56 : wt_actv_nz_out_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1326 = wt_sd_nz_0_57 ? wt_sd_data_0_57 : wt_actv_data_out_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1327 = _T_50633 ? wt_sd_nz_0_57 : wt_actv_nz_out_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1329 = wt_sd_nz_0_58 ? wt_sd_data_0_58 : wt_actv_data_out_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1330 = _T_50633 ? wt_sd_nz_0_58 : wt_actv_nz_out_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1332 = wt_sd_nz_0_59 ? wt_sd_data_0_59 : wt_actv_data_out_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1333 = _T_50633 ? wt_sd_nz_0_59 : wt_actv_nz_out_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1335 = wt_sd_nz_0_60 ? wt_sd_data_0_60 : wt_actv_data_out_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1336 = _T_50633 ? wt_sd_nz_0_60 : wt_actv_nz_out_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1338 = wt_sd_nz_0_61 ? wt_sd_data_0_61 : wt_actv_data_out_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1339 = _T_50633 ? wt_sd_nz_0_61 : wt_actv_nz_out_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1341 = wt_sd_nz_0_62 ? wt_sd_data_0_62 : wt_actv_data_out_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1342 = _T_50633 ? wt_sd_nz_0_62 : wt_actv_nz_out_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1344 = wt_sd_nz_0_63 ? wt_sd_data_0_63 : wt_actv_data_out_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1345 = _T_50633 ? wt_sd_nz_0_63 : wt_actv_nz_out_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1347 = wt_sd_nz_0_64 ? wt_sd_data_0_64 : wt_actv_data_out_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1348 = _T_50633 ? wt_sd_nz_0_64 : wt_actv_nz_out_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1350 = wt_sd_nz_0_65 ? wt_sd_data_0_65 : wt_actv_data_out_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1351 = _T_50633 ? wt_sd_nz_0_65 : wt_actv_nz_out_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1353 = wt_sd_nz_0_66 ? wt_sd_data_0_66 : wt_actv_data_out_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1354 = _T_50633 ? wt_sd_nz_0_66 : wt_actv_nz_out_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1356 = wt_sd_nz_0_67 ? wt_sd_data_0_67 : wt_actv_data_out_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1357 = _T_50633 ? wt_sd_nz_0_67 : wt_actv_nz_out_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1359 = wt_sd_nz_0_68 ? wt_sd_data_0_68 : wt_actv_data_out_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1360 = _T_50633 ? wt_sd_nz_0_68 : wt_actv_nz_out_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1362 = wt_sd_nz_0_69 ? wt_sd_data_0_69 : wt_actv_data_out_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1363 = _T_50633 ? wt_sd_nz_0_69 : wt_actv_nz_out_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1365 = wt_sd_nz_0_70 ? wt_sd_data_0_70 : wt_actv_data_out_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1366 = _T_50633 ? wt_sd_nz_0_70 : wt_actv_nz_out_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1368 = wt_sd_nz_0_71 ? wt_sd_data_0_71 : wt_actv_data_out_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1369 = _T_50633 ? wt_sd_nz_0_71 : wt_actv_nz_out_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1371 = wt_sd_nz_0_72 ? wt_sd_data_0_72 : wt_actv_data_out_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1372 = _T_50633 ? wt_sd_nz_0_72 : wt_actv_nz_out_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1374 = wt_sd_nz_0_73 ? wt_sd_data_0_73 : wt_actv_data_out_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1375 = _T_50633 ? wt_sd_nz_0_73 : wt_actv_nz_out_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1377 = wt_sd_nz_0_74 ? wt_sd_data_0_74 : wt_actv_data_out_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1378 = _T_50633 ? wt_sd_nz_0_74 : wt_actv_nz_out_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1380 = wt_sd_nz_0_75 ? wt_sd_data_0_75 : wt_actv_data_out_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1381 = _T_50633 ? wt_sd_nz_0_75 : wt_actv_nz_out_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1383 = wt_sd_nz_0_76 ? wt_sd_data_0_76 : wt_actv_data_out_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1384 = _T_50633 ? wt_sd_nz_0_76 : wt_actv_nz_out_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1386 = wt_sd_nz_0_77 ? wt_sd_data_0_77 : wt_actv_data_out_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1387 = _T_50633 ? wt_sd_nz_0_77 : wt_actv_nz_out_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1389 = wt_sd_nz_0_78 ? wt_sd_data_0_78 : wt_actv_data_out_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1390 = _T_50633 ? wt_sd_nz_0_78 : wt_actv_nz_out_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1392 = wt_sd_nz_0_79 ? wt_sd_data_0_79 : wt_actv_data_out_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1393 = _T_50633 ? wt_sd_nz_0_79 : wt_actv_nz_out_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1395 = wt_sd_nz_0_80 ? wt_sd_data_0_80 : wt_actv_data_out_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1396 = _T_50633 ? wt_sd_nz_0_80 : wt_actv_nz_out_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1398 = wt_sd_nz_0_81 ? wt_sd_data_0_81 : wt_actv_data_out_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1399 = _T_50633 ? wt_sd_nz_0_81 : wt_actv_nz_out_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1401 = wt_sd_nz_0_82 ? wt_sd_data_0_82 : wt_actv_data_out_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1402 = _T_50633 ? wt_sd_nz_0_82 : wt_actv_nz_out_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1404 = wt_sd_nz_0_83 ? wt_sd_data_0_83 : wt_actv_data_out_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1405 = _T_50633 ? wt_sd_nz_0_83 : wt_actv_nz_out_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1407 = wt_sd_nz_0_84 ? wt_sd_data_0_84 : wt_actv_data_out_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1408 = _T_50633 ? wt_sd_nz_0_84 : wt_actv_nz_out_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1410 = wt_sd_nz_0_85 ? wt_sd_data_0_85 : wt_actv_data_out_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1411 = _T_50633 ? wt_sd_nz_0_85 : wt_actv_nz_out_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1413 = wt_sd_nz_0_86 ? wt_sd_data_0_86 : wt_actv_data_out_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1414 = _T_50633 ? wt_sd_nz_0_86 : wt_actv_nz_out_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1416 = wt_sd_nz_0_87 ? wt_sd_data_0_87 : wt_actv_data_out_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1417 = _T_50633 ? wt_sd_nz_0_87 : wt_actv_nz_out_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1419 = wt_sd_nz_0_88 ? wt_sd_data_0_88 : wt_actv_data_out_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1420 = _T_50633 ? wt_sd_nz_0_88 : wt_actv_nz_out_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1422 = wt_sd_nz_0_89 ? wt_sd_data_0_89 : wt_actv_data_out_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1423 = _T_50633 ? wt_sd_nz_0_89 : wt_actv_nz_out_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1425 = wt_sd_nz_0_90 ? wt_sd_data_0_90 : wt_actv_data_out_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1426 = _T_50633 ? wt_sd_nz_0_90 : wt_actv_nz_out_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1428 = wt_sd_nz_0_91 ? wt_sd_data_0_91 : wt_actv_data_out_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1429 = _T_50633 ? wt_sd_nz_0_91 : wt_actv_nz_out_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1431 = wt_sd_nz_0_92 ? wt_sd_data_0_92 : wt_actv_data_out_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1432 = _T_50633 ? wt_sd_nz_0_92 : wt_actv_nz_out_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1434 = wt_sd_nz_0_93 ? wt_sd_data_0_93 : wt_actv_data_out_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1435 = _T_50633 ? wt_sd_nz_0_93 : wt_actv_nz_out_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1437 = wt_sd_nz_0_94 ? wt_sd_data_0_94 : wt_actv_data_out_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1438 = _T_50633 ? wt_sd_nz_0_94 : wt_actv_nz_out_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1440 = wt_sd_nz_0_95 ? wt_sd_data_0_95 : wt_actv_data_out_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1441 = _T_50633 ? wt_sd_nz_0_95 : wt_actv_nz_out_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1443 = wt_sd_nz_0_96 ? wt_sd_data_0_96 : wt_actv_data_out_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1444 = _T_50633 ? wt_sd_nz_0_96 : wt_actv_nz_out_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1446 = wt_sd_nz_0_97 ? wt_sd_data_0_97 : wt_actv_data_out_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1447 = _T_50633 ? wt_sd_nz_0_97 : wt_actv_nz_out_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1449 = wt_sd_nz_0_98 ? wt_sd_data_0_98 : wt_actv_data_out_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1450 = _T_50633 ? wt_sd_nz_0_98 : wt_actv_nz_out_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1452 = wt_sd_nz_0_99 ? wt_sd_data_0_99 : wt_actv_data_out_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1453 = _T_50633 ? wt_sd_nz_0_99 : wt_actv_nz_out_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1455 = wt_sd_nz_0_100 ? wt_sd_data_0_100 : wt_actv_data_out_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1456 = _T_50633 ? wt_sd_nz_0_100 : wt_actv_nz_out_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1458 = wt_sd_nz_0_101 ? wt_sd_data_0_101 : wt_actv_data_out_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1459 = _T_50633 ? wt_sd_nz_0_101 : wt_actv_nz_out_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1461 = wt_sd_nz_0_102 ? wt_sd_data_0_102 : wt_actv_data_out_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1462 = _T_50633 ? wt_sd_nz_0_102 : wt_actv_nz_out_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1464 = wt_sd_nz_0_103 ? wt_sd_data_0_103 : wt_actv_data_out_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1465 = _T_50633 ? wt_sd_nz_0_103 : wt_actv_nz_out_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1467 = wt_sd_nz_0_104 ? wt_sd_data_0_104 : wt_actv_data_out_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1468 = _T_50633 ? wt_sd_nz_0_104 : wt_actv_nz_out_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1470 = wt_sd_nz_0_105 ? wt_sd_data_0_105 : wt_actv_data_out_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1471 = _T_50633 ? wt_sd_nz_0_105 : wt_actv_nz_out_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1473 = wt_sd_nz_0_106 ? wt_sd_data_0_106 : wt_actv_data_out_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1474 = _T_50633 ? wt_sd_nz_0_106 : wt_actv_nz_out_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1476 = wt_sd_nz_0_107 ? wt_sd_data_0_107 : wt_actv_data_out_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1477 = _T_50633 ? wt_sd_nz_0_107 : wt_actv_nz_out_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1479 = wt_sd_nz_0_108 ? wt_sd_data_0_108 : wt_actv_data_out_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1480 = _T_50633 ? wt_sd_nz_0_108 : wt_actv_nz_out_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1482 = wt_sd_nz_0_109 ? wt_sd_data_0_109 : wt_actv_data_out_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1483 = _T_50633 ? wt_sd_nz_0_109 : wt_actv_nz_out_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1485 = wt_sd_nz_0_110 ? wt_sd_data_0_110 : wt_actv_data_out_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1486 = _T_50633 ? wt_sd_nz_0_110 : wt_actv_nz_out_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1488 = wt_sd_nz_0_111 ? wt_sd_data_0_111 : wt_actv_data_out_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1489 = _T_50633 ? wt_sd_nz_0_111 : wt_actv_nz_out_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1491 = wt_sd_nz_0_112 ? wt_sd_data_0_112 : wt_actv_data_out_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1492 = _T_50633 ? wt_sd_nz_0_112 : wt_actv_nz_out_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1494 = wt_sd_nz_0_113 ? wt_sd_data_0_113 : wt_actv_data_out_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1495 = _T_50633 ? wt_sd_nz_0_113 : wt_actv_nz_out_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1497 = wt_sd_nz_0_114 ? wt_sd_data_0_114 : wt_actv_data_out_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1498 = _T_50633 ? wt_sd_nz_0_114 : wt_actv_nz_out_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1500 = wt_sd_nz_0_115 ? wt_sd_data_0_115 : wt_actv_data_out_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1501 = _T_50633 ? wt_sd_nz_0_115 : wt_actv_nz_out_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1503 = wt_sd_nz_0_116 ? wt_sd_data_0_116 : wt_actv_data_out_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1504 = _T_50633 ? wt_sd_nz_0_116 : wt_actv_nz_out_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1506 = wt_sd_nz_0_117 ? wt_sd_data_0_117 : wt_actv_data_out_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1507 = _T_50633 ? wt_sd_nz_0_117 : wt_actv_nz_out_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1509 = wt_sd_nz_0_118 ? wt_sd_data_0_118 : wt_actv_data_out_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1510 = _T_50633 ? wt_sd_nz_0_118 : wt_actv_nz_out_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1512 = wt_sd_nz_0_119 ? wt_sd_data_0_119 : wt_actv_data_out_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1513 = _T_50633 ? wt_sd_nz_0_119 : wt_actv_nz_out_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1515 = wt_sd_nz_0_120 ? wt_sd_data_0_120 : wt_actv_data_out_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1516 = _T_50633 ? wt_sd_nz_0_120 : wt_actv_nz_out_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1518 = wt_sd_nz_0_121 ? wt_sd_data_0_121 : wt_actv_data_out_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1519 = _T_50633 ? wt_sd_nz_0_121 : wt_actv_nz_out_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1521 = wt_sd_nz_0_122 ? wt_sd_data_0_122 : wt_actv_data_out_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1522 = _T_50633 ? wt_sd_nz_0_122 : wt_actv_nz_out_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1524 = wt_sd_nz_0_123 ? wt_sd_data_0_123 : wt_actv_data_out_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1525 = _T_50633 ? wt_sd_nz_0_123 : wt_actv_nz_out_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1527 = wt_sd_nz_0_124 ? wt_sd_data_0_124 : wt_actv_data_out_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1528 = _T_50633 ? wt_sd_nz_0_124 : wt_actv_nz_out_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1530 = wt_sd_nz_0_125 ? wt_sd_data_0_125 : wt_actv_data_out_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1531 = _T_50633 ? wt_sd_nz_0_125 : wt_actv_nz_out_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1533 = wt_sd_nz_0_126 ? wt_sd_data_0_126 : wt_actv_data_out_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1534 = _T_50633 ? wt_sd_nz_0_126 : wt_actv_nz_out_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1536 = wt_sd_nz_0_127 ? wt_sd_data_0_127 : wt_actv_data_out_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 147:37]
  assign _GEN_1537 = _T_50633 ? wt_sd_nz_0_127 : wt_actv_nz_out_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 145:61]
  assign _GEN_1539 = dat_pre_pvld ? dat_pre_nz_0 : dat_actv_nz_reg_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1540 = dat_pre_pvld ? dat_pre_nz_1 : dat_actv_nz_reg_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1541 = dat_pre_pvld ? dat_pre_nz_2 : dat_actv_nz_reg_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1542 = dat_pre_pvld ? dat_pre_nz_3 : dat_actv_nz_reg_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1543 = dat_pre_pvld ? dat_pre_nz_4 : dat_actv_nz_reg_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1544 = dat_pre_pvld ? dat_pre_nz_5 : dat_actv_nz_reg_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1545 = dat_pre_pvld ? dat_pre_nz_6 : dat_actv_nz_reg_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1546 = dat_pre_pvld ? dat_pre_nz_7 : dat_actv_nz_reg_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1547 = dat_pre_pvld ? dat_pre_nz_8 : dat_actv_nz_reg_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1548 = dat_pre_pvld ? dat_pre_nz_9 : dat_actv_nz_reg_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1549 = dat_pre_pvld ? dat_pre_nz_10 : dat_actv_nz_reg_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1550 = dat_pre_pvld ? dat_pre_nz_11 : dat_actv_nz_reg_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1551 = dat_pre_pvld ? dat_pre_nz_12 : dat_actv_nz_reg_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1552 = dat_pre_pvld ? dat_pre_nz_13 : dat_actv_nz_reg_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1553 = dat_pre_pvld ? dat_pre_nz_14 : dat_actv_nz_reg_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1554 = dat_pre_pvld ? dat_pre_nz_15 : dat_actv_nz_reg_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1555 = dat_pre_pvld ? dat_pre_nz_16 : dat_actv_nz_reg_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1556 = dat_pre_pvld ? dat_pre_nz_17 : dat_actv_nz_reg_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1557 = dat_pre_pvld ? dat_pre_nz_18 : dat_actv_nz_reg_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1558 = dat_pre_pvld ? dat_pre_nz_19 : dat_actv_nz_reg_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1559 = dat_pre_pvld ? dat_pre_nz_20 : dat_actv_nz_reg_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1560 = dat_pre_pvld ? dat_pre_nz_21 : dat_actv_nz_reg_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1561 = dat_pre_pvld ? dat_pre_nz_22 : dat_actv_nz_reg_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1562 = dat_pre_pvld ? dat_pre_nz_23 : dat_actv_nz_reg_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1563 = dat_pre_pvld ? dat_pre_nz_24 : dat_actv_nz_reg_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1564 = dat_pre_pvld ? dat_pre_nz_25 : dat_actv_nz_reg_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1565 = dat_pre_pvld ? dat_pre_nz_26 : dat_actv_nz_reg_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1566 = dat_pre_pvld ? dat_pre_nz_27 : dat_actv_nz_reg_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1567 = dat_pre_pvld ? dat_pre_nz_28 : dat_actv_nz_reg_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1568 = dat_pre_pvld ? dat_pre_nz_29 : dat_actv_nz_reg_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1569 = dat_pre_pvld ? dat_pre_nz_30 : dat_actv_nz_reg_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1570 = dat_pre_pvld ? dat_pre_nz_31 : dat_actv_nz_reg_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1571 = dat_pre_pvld ? dat_pre_nz_32 : dat_actv_nz_reg_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1572 = dat_pre_pvld ? dat_pre_nz_33 : dat_actv_nz_reg_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1573 = dat_pre_pvld ? dat_pre_nz_34 : dat_actv_nz_reg_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1574 = dat_pre_pvld ? dat_pre_nz_35 : dat_actv_nz_reg_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1575 = dat_pre_pvld ? dat_pre_nz_36 : dat_actv_nz_reg_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1576 = dat_pre_pvld ? dat_pre_nz_37 : dat_actv_nz_reg_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1577 = dat_pre_pvld ? dat_pre_nz_38 : dat_actv_nz_reg_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1578 = dat_pre_pvld ? dat_pre_nz_39 : dat_actv_nz_reg_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1579 = dat_pre_pvld ? dat_pre_nz_40 : dat_actv_nz_reg_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1580 = dat_pre_pvld ? dat_pre_nz_41 : dat_actv_nz_reg_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1581 = dat_pre_pvld ? dat_pre_nz_42 : dat_actv_nz_reg_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1582 = dat_pre_pvld ? dat_pre_nz_43 : dat_actv_nz_reg_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1583 = dat_pre_pvld ? dat_pre_nz_44 : dat_actv_nz_reg_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1584 = dat_pre_pvld ? dat_pre_nz_45 : dat_actv_nz_reg_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1585 = dat_pre_pvld ? dat_pre_nz_46 : dat_actv_nz_reg_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1586 = dat_pre_pvld ? dat_pre_nz_47 : dat_actv_nz_reg_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1587 = dat_pre_pvld ? dat_pre_nz_48 : dat_actv_nz_reg_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1588 = dat_pre_pvld ? dat_pre_nz_49 : dat_actv_nz_reg_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1589 = dat_pre_pvld ? dat_pre_nz_50 : dat_actv_nz_reg_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1590 = dat_pre_pvld ? dat_pre_nz_51 : dat_actv_nz_reg_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1591 = dat_pre_pvld ? dat_pre_nz_52 : dat_actv_nz_reg_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1592 = dat_pre_pvld ? dat_pre_nz_53 : dat_actv_nz_reg_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1593 = dat_pre_pvld ? dat_pre_nz_54 : dat_actv_nz_reg_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1594 = dat_pre_pvld ? dat_pre_nz_55 : dat_actv_nz_reg_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1595 = dat_pre_pvld ? dat_pre_nz_56 : dat_actv_nz_reg_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1596 = dat_pre_pvld ? dat_pre_nz_57 : dat_actv_nz_reg_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1597 = dat_pre_pvld ? dat_pre_nz_58 : dat_actv_nz_reg_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1598 = dat_pre_pvld ? dat_pre_nz_59 : dat_actv_nz_reg_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1599 = dat_pre_pvld ? dat_pre_nz_60 : dat_actv_nz_reg_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1600 = dat_pre_pvld ? dat_pre_nz_61 : dat_actv_nz_reg_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1601 = dat_pre_pvld ? dat_pre_nz_62 : dat_actv_nz_reg_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1602 = dat_pre_pvld ? dat_pre_nz_63 : dat_actv_nz_reg_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1603 = dat_pre_pvld ? dat_pre_nz_64 : dat_actv_nz_reg_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1604 = dat_pre_pvld ? dat_pre_nz_65 : dat_actv_nz_reg_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1605 = dat_pre_pvld ? dat_pre_nz_66 : dat_actv_nz_reg_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1606 = dat_pre_pvld ? dat_pre_nz_67 : dat_actv_nz_reg_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1607 = dat_pre_pvld ? dat_pre_nz_68 : dat_actv_nz_reg_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1608 = dat_pre_pvld ? dat_pre_nz_69 : dat_actv_nz_reg_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1609 = dat_pre_pvld ? dat_pre_nz_70 : dat_actv_nz_reg_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1610 = dat_pre_pvld ? dat_pre_nz_71 : dat_actv_nz_reg_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1611 = dat_pre_pvld ? dat_pre_nz_72 : dat_actv_nz_reg_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1612 = dat_pre_pvld ? dat_pre_nz_73 : dat_actv_nz_reg_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1613 = dat_pre_pvld ? dat_pre_nz_74 : dat_actv_nz_reg_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1614 = dat_pre_pvld ? dat_pre_nz_75 : dat_actv_nz_reg_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1615 = dat_pre_pvld ? dat_pre_nz_76 : dat_actv_nz_reg_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1616 = dat_pre_pvld ? dat_pre_nz_77 : dat_actv_nz_reg_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1617 = dat_pre_pvld ? dat_pre_nz_78 : dat_actv_nz_reg_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1618 = dat_pre_pvld ? dat_pre_nz_79 : dat_actv_nz_reg_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1619 = dat_pre_pvld ? dat_pre_nz_80 : dat_actv_nz_reg_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1620 = dat_pre_pvld ? dat_pre_nz_81 : dat_actv_nz_reg_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1621 = dat_pre_pvld ? dat_pre_nz_82 : dat_actv_nz_reg_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1622 = dat_pre_pvld ? dat_pre_nz_83 : dat_actv_nz_reg_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1623 = dat_pre_pvld ? dat_pre_nz_84 : dat_actv_nz_reg_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1624 = dat_pre_pvld ? dat_pre_nz_85 : dat_actv_nz_reg_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1625 = dat_pre_pvld ? dat_pre_nz_86 : dat_actv_nz_reg_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1626 = dat_pre_pvld ? dat_pre_nz_87 : dat_actv_nz_reg_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1627 = dat_pre_pvld ? dat_pre_nz_88 : dat_actv_nz_reg_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1628 = dat_pre_pvld ? dat_pre_nz_89 : dat_actv_nz_reg_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1629 = dat_pre_pvld ? dat_pre_nz_90 : dat_actv_nz_reg_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1630 = dat_pre_pvld ? dat_pre_nz_91 : dat_actv_nz_reg_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1631 = dat_pre_pvld ? dat_pre_nz_92 : dat_actv_nz_reg_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1632 = dat_pre_pvld ? dat_pre_nz_93 : dat_actv_nz_reg_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1633 = dat_pre_pvld ? dat_pre_nz_94 : dat_actv_nz_reg_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1634 = dat_pre_pvld ? dat_pre_nz_95 : dat_actv_nz_reg_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1635 = dat_pre_pvld ? dat_pre_nz_96 : dat_actv_nz_reg_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1636 = dat_pre_pvld ? dat_pre_nz_97 : dat_actv_nz_reg_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1637 = dat_pre_pvld ? dat_pre_nz_98 : dat_actv_nz_reg_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1638 = dat_pre_pvld ? dat_pre_nz_99 : dat_actv_nz_reg_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1639 = dat_pre_pvld ? dat_pre_nz_100 : dat_actv_nz_reg_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1640 = dat_pre_pvld ? dat_pre_nz_101 : dat_actv_nz_reg_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1641 = dat_pre_pvld ? dat_pre_nz_102 : dat_actv_nz_reg_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1642 = dat_pre_pvld ? dat_pre_nz_103 : dat_actv_nz_reg_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1643 = dat_pre_pvld ? dat_pre_nz_104 : dat_actv_nz_reg_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1644 = dat_pre_pvld ? dat_pre_nz_105 : dat_actv_nz_reg_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1645 = dat_pre_pvld ? dat_pre_nz_106 : dat_actv_nz_reg_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1646 = dat_pre_pvld ? dat_pre_nz_107 : dat_actv_nz_reg_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1647 = dat_pre_pvld ? dat_pre_nz_108 : dat_actv_nz_reg_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1648 = dat_pre_pvld ? dat_pre_nz_109 : dat_actv_nz_reg_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1649 = dat_pre_pvld ? dat_pre_nz_110 : dat_actv_nz_reg_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1650 = dat_pre_pvld ? dat_pre_nz_111 : dat_actv_nz_reg_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1651 = dat_pre_pvld ? dat_pre_nz_112 : dat_actv_nz_reg_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1652 = dat_pre_pvld ? dat_pre_nz_113 : dat_actv_nz_reg_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1653 = dat_pre_pvld ? dat_pre_nz_114 : dat_actv_nz_reg_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1654 = dat_pre_pvld ? dat_pre_nz_115 : dat_actv_nz_reg_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1655 = dat_pre_pvld ? dat_pre_nz_116 : dat_actv_nz_reg_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1656 = dat_pre_pvld ? dat_pre_nz_117 : dat_actv_nz_reg_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1657 = dat_pre_pvld ? dat_pre_nz_118 : dat_actv_nz_reg_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1658 = dat_pre_pvld ? dat_pre_nz_119 : dat_actv_nz_reg_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1659 = dat_pre_pvld ? dat_pre_nz_120 : dat_actv_nz_reg_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1660 = dat_pre_pvld ? dat_pre_nz_121 : dat_actv_nz_reg_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1661 = dat_pre_pvld ? dat_pre_nz_122 : dat_actv_nz_reg_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1662 = dat_pre_pvld ? dat_pre_nz_123 : dat_actv_nz_reg_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1663 = dat_pre_pvld ? dat_pre_nz_124 : dat_actv_nz_reg_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1664 = dat_pre_pvld ? dat_pre_nz_125 : dat_actv_nz_reg_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1665 = dat_pre_pvld ? dat_pre_nz_126 : dat_actv_nz_reg_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _GEN_1666 = dat_pre_pvld ? dat_pre_nz_127 : dat_actv_nz_reg_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 167:27]
  assign _T_73569 = dat_pre_pvld & dat_pre_nz_0; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73570 = dat_pre_pvld & dat_pre_nz_1; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73571 = dat_pre_pvld & dat_pre_nz_2; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73572 = dat_pre_pvld & dat_pre_nz_3; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73573 = dat_pre_pvld & dat_pre_nz_4; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73574 = dat_pre_pvld & dat_pre_nz_5; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73575 = dat_pre_pvld & dat_pre_nz_6; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73576 = dat_pre_pvld & dat_pre_nz_7; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73577 = dat_pre_pvld & dat_pre_nz_8; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73578 = dat_pre_pvld & dat_pre_nz_9; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73579 = dat_pre_pvld & dat_pre_nz_10; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73580 = dat_pre_pvld & dat_pre_nz_11; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73581 = dat_pre_pvld & dat_pre_nz_12; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73582 = dat_pre_pvld & dat_pre_nz_13; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73583 = dat_pre_pvld & dat_pre_nz_14; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73584 = dat_pre_pvld & dat_pre_nz_15; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73585 = dat_pre_pvld & dat_pre_nz_16; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73586 = dat_pre_pvld & dat_pre_nz_17; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73587 = dat_pre_pvld & dat_pre_nz_18; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73588 = dat_pre_pvld & dat_pre_nz_19; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73589 = dat_pre_pvld & dat_pre_nz_20; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73590 = dat_pre_pvld & dat_pre_nz_21; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73591 = dat_pre_pvld & dat_pre_nz_22; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73592 = dat_pre_pvld & dat_pre_nz_23; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73593 = dat_pre_pvld & dat_pre_nz_24; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73594 = dat_pre_pvld & dat_pre_nz_25; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73595 = dat_pre_pvld & dat_pre_nz_26; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73596 = dat_pre_pvld & dat_pre_nz_27; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73597 = dat_pre_pvld & dat_pre_nz_28; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73598 = dat_pre_pvld & dat_pre_nz_29; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73599 = dat_pre_pvld & dat_pre_nz_30; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73600 = dat_pre_pvld & dat_pre_nz_31; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73601 = dat_pre_pvld & dat_pre_nz_32; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73602 = dat_pre_pvld & dat_pre_nz_33; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73603 = dat_pre_pvld & dat_pre_nz_34; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73604 = dat_pre_pvld & dat_pre_nz_35; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73605 = dat_pre_pvld & dat_pre_nz_36; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73606 = dat_pre_pvld & dat_pre_nz_37; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73607 = dat_pre_pvld & dat_pre_nz_38; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73608 = dat_pre_pvld & dat_pre_nz_39; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73609 = dat_pre_pvld & dat_pre_nz_40; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73610 = dat_pre_pvld & dat_pre_nz_41; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73611 = dat_pre_pvld & dat_pre_nz_42; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73612 = dat_pre_pvld & dat_pre_nz_43; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73613 = dat_pre_pvld & dat_pre_nz_44; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73614 = dat_pre_pvld & dat_pre_nz_45; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73615 = dat_pre_pvld & dat_pre_nz_46; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73616 = dat_pre_pvld & dat_pre_nz_47; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73617 = dat_pre_pvld & dat_pre_nz_48; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73618 = dat_pre_pvld & dat_pre_nz_49; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73619 = dat_pre_pvld & dat_pre_nz_50; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73620 = dat_pre_pvld & dat_pre_nz_51; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73621 = dat_pre_pvld & dat_pre_nz_52; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73622 = dat_pre_pvld & dat_pre_nz_53; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73623 = dat_pre_pvld & dat_pre_nz_54; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73624 = dat_pre_pvld & dat_pre_nz_55; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73625 = dat_pre_pvld & dat_pre_nz_56; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73626 = dat_pre_pvld & dat_pre_nz_57; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73627 = dat_pre_pvld & dat_pre_nz_58; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73628 = dat_pre_pvld & dat_pre_nz_59; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73629 = dat_pre_pvld & dat_pre_nz_60; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73630 = dat_pre_pvld & dat_pre_nz_61; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73631 = dat_pre_pvld & dat_pre_nz_62; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73632 = dat_pre_pvld & dat_pre_nz_63; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73633 = dat_pre_pvld & dat_pre_nz_64; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73634 = dat_pre_pvld & dat_pre_nz_65; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73635 = dat_pre_pvld & dat_pre_nz_66; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73636 = dat_pre_pvld & dat_pre_nz_67; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73637 = dat_pre_pvld & dat_pre_nz_68; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73638 = dat_pre_pvld & dat_pre_nz_69; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73639 = dat_pre_pvld & dat_pre_nz_70; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73640 = dat_pre_pvld & dat_pre_nz_71; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73641 = dat_pre_pvld & dat_pre_nz_72; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73642 = dat_pre_pvld & dat_pre_nz_73; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73643 = dat_pre_pvld & dat_pre_nz_74; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73644 = dat_pre_pvld & dat_pre_nz_75; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73645 = dat_pre_pvld & dat_pre_nz_76; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73646 = dat_pre_pvld & dat_pre_nz_77; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73647 = dat_pre_pvld & dat_pre_nz_78; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73648 = dat_pre_pvld & dat_pre_nz_79; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73649 = dat_pre_pvld & dat_pre_nz_80; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73650 = dat_pre_pvld & dat_pre_nz_81; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73651 = dat_pre_pvld & dat_pre_nz_82; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73652 = dat_pre_pvld & dat_pre_nz_83; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73653 = dat_pre_pvld & dat_pre_nz_84; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73654 = dat_pre_pvld & dat_pre_nz_85; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73655 = dat_pre_pvld & dat_pre_nz_86; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73656 = dat_pre_pvld & dat_pre_nz_87; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73657 = dat_pre_pvld & dat_pre_nz_88; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73658 = dat_pre_pvld & dat_pre_nz_89; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73659 = dat_pre_pvld & dat_pre_nz_90; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73660 = dat_pre_pvld & dat_pre_nz_91; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73661 = dat_pre_pvld & dat_pre_nz_92; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73662 = dat_pre_pvld & dat_pre_nz_93; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73663 = dat_pre_pvld & dat_pre_nz_94; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73664 = dat_pre_pvld & dat_pre_nz_95; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73665 = dat_pre_pvld & dat_pre_nz_96; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73666 = dat_pre_pvld & dat_pre_nz_97; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73667 = dat_pre_pvld & dat_pre_nz_98; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73668 = dat_pre_pvld & dat_pre_nz_99; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73669 = dat_pre_pvld & dat_pre_nz_100; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73670 = dat_pre_pvld & dat_pre_nz_101; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73671 = dat_pre_pvld & dat_pre_nz_102; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73672 = dat_pre_pvld & dat_pre_nz_103; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73673 = dat_pre_pvld & dat_pre_nz_104; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73674 = dat_pre_pvld & dat_pre_nz_105; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73675 = dat_pre_pvld & dat_pre_nz_106; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73676 = dat_pre_pvld & dat_pre_nz_107; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73677 = dat_pre_pvld & dat_pre_nz_108; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73678 = dat_pre_pvld & dat_pre_nz_109; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73679 = dat_pre_pvld & dat_pre_nz_110; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73680 = dat_pre_pvld & dat_pre_nz_111; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73681 = dat_pre_pvld & dat_pre_nz_112; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73682 = dat_pre_pvld & dat_pre_nz_113; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73683 = dat_pre_pvld & dat_pre_nz_114; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73684 = dat_pre_pvld & dat_pre_nz_115; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73685 = dat_pre_pvld & dat_pre_nz_116; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73686 = dat_pre_pvld & dat_pre_nz_117; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73687 = dat_pre_pvld & dat_pre_nz_118; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73688 = dat_pre_pvld & dat_pre_nz_119; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73689 = dat_pre_pvld & dat_pre_nz_120; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73690 = dat_pre_pvld & dat_pre_nz_121; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73691 = dat_pre_pvld & dat_pre_nz_122; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73692 = dat_pre_pvld & dat_pre_nz_123; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73693 = dat_pre_pvld & dat_pre_nz_124; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73694 = dat_pre_pvld & dat_pre_nz_125; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73695 = dat_pre_pvld & dat_pre_nz_126; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign _T_73696 = dat_pre_pvld & dat_pre_nz_127; // @[NV_NVDLA_CMAC_CORE_active.scala 171:30]
  assign io_dat_actv_data_0_0 = dat_actv_data_reg_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_1 = dat_actv_data_reg_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_2 = dat_actv_data_reg_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_3 = dat_actv_data_reg_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_4 = dat_actv_data_reg_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_5 = dat_actv_data_reg_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_6 = dat_actv_data_reg_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_7 = dat_actv_data_reg_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_8 = dat_actv_data_reg_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_9 = dat_actv_data_reg_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_10 = dat_actv_data_reg_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_11 = dat_actv_data_reg_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_12 = dat_actv_data_reg_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_13 = dat_actv_data_reg_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_14 = dat_actv_data_reg_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_15 = dat_actv_data_reg_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_16 = dat_actv_data_reg_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_17 = dat_actv_data_reg_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_18 = dat_actv_data_reg_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_19 = dat_actv_data_reg_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_20 = dat_actv_data_reg_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_21 = dat_actv_data_reg_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_22 = dat_actv_data_reg_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_23 = dat_actv_data_reg_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_24 = dat_actv_data_reg_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_25 = dat_actv_data_reg_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_26 = dat_actv_data_reg_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_27 = dat_actv_data_reg_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_28 = dat_actv_data_reg_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_29 = dat_actv_data_reg_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_30 = dat_actv_data_reg_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_31 = dat_actv_data_reg_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_32 = dat_actv_data_reg_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_33 = dat_actv_data_reg_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_34 = dat_actv_data_reg_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_35 = dat_actv_data_reg_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_36 = dat_actv_data_reg_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_37 = dat_actv_data_reg_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_38 = dat_actv_data_reg_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_39 = dat_actv_data_reg_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_40 = dat_actv_data_reg_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_41 = dat_actv_data_reg_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_42 = dat_actv_data_reg_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_43 = dat_actv_data_reg_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_44 = dat_actv_data_reg_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_45 = dat_actv_data_reg_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_46 = dat_actv_data_reg_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_47 = dat_actv_data_reg_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_48 = dat_actv_data_reg_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_49 = dat_actv_data_reg_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_50 = dat_actv_data_reg_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_51 = dat_actv_data_reg_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_52 = dat_actv_data_reg_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_53 = dat_actv_data_reg_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_54 = dat_actv_data_reg_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_55 = dat_actv_data_reg_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_56 = dat_actv_data_reg_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_57 = dat_actv_data_reg_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_58 = dat_actv_data_reg_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_59 = dat_actv_data_reg_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_60 = dat_actv_data_reg_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_61 = dat_actv_data_reg_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_62 = dat_actv_data_reg_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_63 = dat_actv_data_reg_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_64 = dat_actv_data_reg_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_65 = dat_actv_data_reg_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_66 = dat_actv_data_reg_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_67 = dat_actv_data_reg_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_68 = dat_actv_data_reg_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_69 = dat_actv_data_reg_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_70 = dat_actv_data_reg_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_71 = dat_actv_data_reg_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_72 = dat_actv_data_reg_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_73 = dat_actv_data_reg_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_74 = dat_actv_data_reg_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_75 = dat_actv_data_reg_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_76 = dat_actv_data_reg_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_77 = dat_actv_data_reg_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_78 = dat_actv_data_reg_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_79 = dat_actv_data_reg_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_80 = dat_actv_data_reg_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_81 = dat_actv_data_reg_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_82 = dat_actv_data_reg_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_83 = dat_actv_data_reg_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_84 = dat_actv_data_reg_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_85 = dat_actv_data_reg_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_86 = dat_actv_data_reg_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_87 = dat_actv_data_reg_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_88 = dat_actv_data_reg_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_89 = dat_actv_data_reg_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_90 = dat_actv_data_reg_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_91 = dat_actv_data_reg_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_92 = dat_actv_data_reg_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_93 = dat_actv_data_reg_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_94 = dat_actv_data_reg_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_95 = dat_actv_data_reg_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_96 = dat_actv_data_reg_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_97 = dat_actv_data_reg_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_98 = dat_actv_data_reg_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_99 = dat_actv_data_reg_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_100 = dat_actv_data_reg_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_101 = dat_actv_data_reg_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_102 = dat_actv_data_reg_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_103 = dat_actv_data_reg_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_104 = dat_actv_data_reg_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_105 = dat_actv_data_reg_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_106 = dat_actv_data_reg_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_107 = dat_actv_data_reg_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_108 = dat_actv_data_reg_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_109 = dat_actv_data_reg_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_110 = dat_actv_data_reg_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_111 = dat_actv_data_reg_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_112 = dat_actv_data_reg_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_113 = dat_actv_data_reg_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_114 = dat_actv_data_reg_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_115 = dat_actv_data_reg_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_116 = dat_actv_data_reg_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_117 = dat_actv_data_reg_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_118 = dat_actv_data_reg_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_119 = dat_actv_data_reg_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_120 = dat_actv_data_reg_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_121 = dat_actv_data_reg_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_122 = dat_actv_data_reg_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_123 = dat_actv_data_reg_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_124 = dat_actv_data_reg_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_125 = dat_actv_data_reg_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_126 = dat_actv_data_reg_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_data_0_127 = dat_actv_data_reg_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 187:22]
  assign io_dat_actv_nz_0_0 = dat_actv_nz_reg_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_1 = dat_actv_nz_reg_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_2 = dat_actv_nz_reg_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_3 = dat_actv_nz_reg_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_4 = dat_actv_nz_reg_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_5 = dat_actv_nz_reg_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_6 = dat_actv_nz_reg_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_7 = dat_actv_nz_reg_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_8 = dat_actv_nz_reg_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_9 = dat_actv_nz_reg_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_10 = dat_actv_nz_reg_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_11 = dat_actv_nz_reg_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_12 = dat_actv_nz_reg_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_13 = dat_actv_nz_reg_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_14 = dat_actv_nz_reg_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_15 = dat_actv_nz_reg_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_16 = dat_actv_nz_reg_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_17 = dat_actv_nz_reg_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_18 = dat_actv_nz_reg_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_19 = dat_actv_nz_reg_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_20 = dat_actv_nz_reg_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_21 = dat_actv_nz_reg_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_22 = dat_actv_nz_reg_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_23 = dat_actv_nz_reg_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_24 = dat_actv_nz_reg_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_25 = dat_actv_nz_reg_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_26 = dat_actv_nz_reg_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_27 = dat_actv_nz_reg_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_28 = dat_actv_nz_reg_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_29 = dat_actv_nz_reg_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_30 = dat_actv_nz_reg_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_31 = dat_actv_nz_reg_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_32 = dat_actv_nz_reg_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_33 = dat_actv_nz_reg_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_34 = dat_actv_nz_reg_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_35 = dat_actv_nz_reg_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_36 = dat_actv_nz_reg_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_37 = dat_actv_nz_reg_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_38 = dat_actv_nz_reg_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_39 = dat_actv_nz_reg_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_40 = dat_actv_nz_reg_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_41 = dat_actv_nz_reg_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_42 = dat_actv_nz_reg_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_43 = dat_actv_nz_reg_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_44 = dat_actv_nz_reg_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_45 = dat_actv_nz_reg_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_46 = dat_actv_nz_reg_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_47 = dat_actv_nz_reg_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_48 = dat_actv_nz_reg_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_49 = dat_actv_nz_reg_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_50 = dat_actv_nz_reg_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_51 = dat_actv_nz_reg_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_52 = dat_actv_nz_reg_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_53 = dat_actv_nz_reg_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_54 = dat_actv_nz_reg_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_55 = dat_actv_nz_reg_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_56 = dat_actv_nz_reg_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_57 = dat_actv_nz_reg_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_58 = dat_actv_nz_reg_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_59 = dat_actv_nz_reg_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_60 = dat_actv_nz_reg_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_61 = dat_actv_nz_reg_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_62 = dat_actv_nz_reg_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_63 = dat_actv_nz_reg_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_64 = dat_actv_nz_reg_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_65 = dat_actv_nz_reg_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_66 = dat_actv_nz_reg_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_67 = dat_actv_nz_reg_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_68 = dat_actv_nz_reg_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_69 = dat_actv_nz_reg_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_70 = dat_actv_nz_reg_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_71 = dat_actv_nz_reg_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_72 = dat_actv_nz_reg_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_73 = dat_actv_nz_reg_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_74 = dat_actv_nz_reg_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_75 = dat_actv_nz_reg_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_76 = dat_actv_nz_reg_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_77 = dat_actv_nz_reg_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_78 = dat_actv_nz_reg_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_79 = dat_actv_nz_reg_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_80 = dat_actv_nz_reg_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_81 = dat_actv_nz_reg_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_82 = dat_actv_nz_reg_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_83 = dat_actv_nz_reg_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_84 = dat_actv_nz_reg_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_85 = dat_actv_nz_reg_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_86 = dat_actv_nz_reg_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_87 = dat_actv_nz_reg_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_88 = dat_actv_nz_reg_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_89 = dat_actv_nz_reg_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_90 = dat_actv_nz_reg_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_91 = dat_actv_nz_reg_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_92 = dat_actv_nz_reg_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_93 = dat_actv_nz_reg_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_94 = dat_actv_nz_reg_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_95 = dat_actv_nz_reg_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_96 = dat_actv_nz_reg_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_97 = dat_actv_nz_reg_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_98 = dat_actv_nz_reg_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_99 = dat_actv_nz_reg_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_100 = dat_actv_nz_reg_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_101 = dat_actv_nz_reg_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_102 = dat_actv_nz_reg_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_103 = dat_actv_nz_reg_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_104 = dat_actv_nz_reg_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_105 = dat_actv_nz_reg_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_106 = dat_actv_nz_reg_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_107 = dat_actv_nz_reg_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_108 = dat_actv_nz_reg_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_109 = dat_actv_nz_reg_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_110 = dat_actv_nz_reg_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_111 = dat_actv_nz_reg_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_112 = dat_actv_nz_reg_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_113 = dat_actv_nz_reg_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_114 = dat_actv_nz_reg_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_115 = dat_actv_nz_reg_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_116 = dat_actv_nz_reg_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_117 = dat_actv_nz_reg_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_118 = dat_actv_nz_reg_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_119 = dat_actv_nz_reg_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_120 = dat_actv_nz_reg_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_121 = dat_actv_nz_reg_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_122 = dat_actv_nz_reg_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_123 = dat_actv_nz_reg_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_124 = dat_actv_nz_reg_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_125 = dat_actv_nz_reg_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_126 = dat_actv_nz_reg_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_nz_0_127 = dat_actv_nz_reg_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 188:20]
  assign io_dat_actv_pvld_0_0 = dat_actv_pvld_reg_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_1 = dat_actv_pvld_reg_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_2 = dat_actv_pvld_reg_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_3 = dat_actv_pvld_reg_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_4 = dat_actv_pvld_reg_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_5 = dat_actv_pvld_reg_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_6 = dat_actv_pvld_reg_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_7 = dat_actv_pvld_reg_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_8 = dat_actv_pvld_reg_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_9 = dat_actv_pvld_reg_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_10 = dat_actv_pvld_reg_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_11 = dat_actv_pvld_reg_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_12 = dat_actv_pvld_reg_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_13 = dat_actv_pvld_reg_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_14 = dat_actv_pvld_reg_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_15 = dat_actv_pvld_reg_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_16 = dat_actv_pvld_reg_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_17 = dat_actv_pvld_reg_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_18 = dat_actv_pvld_reg_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_19 = dat_actv_pvld_reg_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_20 = dat_actv_pvld_reg_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_21 = dat_actv_pvld_reg_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_22 = dat_actv_pvld_reg_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_23 = dat_actv_pvld_reg_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_24 = dat_actv_pvld_reg_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_25 = dat_actv_pvld_reg_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_26 = dat_actv_pvld_reg_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_27 = dat_actv_pvld_reg_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_28 = dat_actv_pvld_reg_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_29 = dat_actv_pvld_reg_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_30 = dat_actv_pvld_reg_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_31 = dat_actv_pvld_reg_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_32 = dat_actv_pvld_reg_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_33 = dat_actv_pvld_reg_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_34 = dat_actv_pvld_reg_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_35 = dat_actv_pvld_reg_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_36 = dat_actv_pvld_reg_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_37 = dat_actv_pvld_reg_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_38 = dat_actv_pvld_reg_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_39 = dat_actv_pvld_reg_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_40 = dat_actv_pvld_reg_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_41 = dat_actv_pvld_reg_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_42 = dat_actv_pvld_reg_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_43 = dat_actv_pvld_reg_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_44 = dat_actv_pvld_reg_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_45 = dat_actv_pvld_reg_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_46 = dat_actv_pvld_reg_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_47 = dat_actv_pvld_reg_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_48 = dat_actv_pvld_reg_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_49 = dat_actv_pvld_reg_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_50 = dat_actv_pvld_reg_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_51 = dat_actv_pvld_reg_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_52 = dat_actv_pvld_reg_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_53 = dat_actv_pvld_reg_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_54 = dat_actv_pvld_reg_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_55 = dat_actv_pvld_reg_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_56 = dat_actv_pvld_reg_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_57 = dat_actv_pvld_reg_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_58 = dat_actv_pvld_reg_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_59 = dat_actv_pvld_reg_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_60 = dat_actv_pvld_reg_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_61 = dat_actv_pvld_reg_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_62 = dat_actv_pvld_reg_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_63 = dat_actv_pvld_reg_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_64 = dat_actv_pvld_reg_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_65 = dat_actv_pvld_reg_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_66 = dat_actv_pvld_reg_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_67 = dat_actv_pvld_reg_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_68 = dat_actv_pvld_reg_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_69 = dat_actv_pvld_reg_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_70 = dat_actv_pvld_reg_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_71 = dat_actv_pvld_reg_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_72 = dat_actv_pvld_reg_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_73 = dat_actv_pvld_reg_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_74 = dat_actv_pvld_reg_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_75 = dat_actv_pvld_reg_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_76 = dat_actv_pvld_reg_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_77 = dat_actv_pvld_reg_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_78 = dat_actv_pvld_reg_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_79 = dat_actv_pvld_reg_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_80 = dat_actv_pvld_reg_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_81 = dat_actv_pvld_reg_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_82 = dat_actv_pvld_reg_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_83 = dat_actv_pvld_reg_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_84 = dat_actv_pvld_reg_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_85 = dat_actv_pvld_reg_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_86 = dat_actv_pvld_reg_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_87 = dat_actv_pvld_reg_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_88 = dat_actv_pvld_reg_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_89 = dat_actv_pvld_reg_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_90 = dat_actv_pvld_reg_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_91 = dat_actv_pvld_reg_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_92 = dat_actv_pvld_reg_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_93 = dat_actv_pvld_reg_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_94 = dat_actv_pvld_reg_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_95 = dat_actv_pvld_reg_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_96 = dat_actv_pvld_reg_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_97 = dat_actv_pvld_reg_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_98 = dat_actv_pvld_reg_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_99 = dat_actv_pvld_reg_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_100 = dat_actv_pvld_reg_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_101 = dat_actv_pvld_reg_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_102 = dat_actv_pvld_reg_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_103 = dat_actv_pvld_reg_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_104 = dat_actv_pvld_reg_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_105 = dat_actv_pvld_reg_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_106 = dat_actv_pvld_reg_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_107 = dat_actv_pvld_reg_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_108 = dat_actv_pvld_reg_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_109 = dat_actv_pvld_reg_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_110 = dat_actv_pvld_reg_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_111 = dat_actv_pvld_reg_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_112 = dat_actv_pvld_reg_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_113 = dat_actv_pvld_reg_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_114 = dat_actv_pvld_reg_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_115 = dat_actv_pvld_reg_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_116 = dat_actv_pvld_reg_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_117 = dat_actv_pvld_reg_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_118 = dat_actv_pvld_reg_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_119 = dat_actv_pvld_reg_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_120 = dat_actv_pvld_reg_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_121 = dat_actv_pvld_reg_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_122 = dat_actv_pvld_reg_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_123 = dat_actv_pvld_reg_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_124 = dat_actv_pvld_reg_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_125 = dat_actv_pvld_reg_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_126 = dat_actv_pvld_reg_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_dat_actv_pvld_0_127 = dat_actv_pvld_reg_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 186:22]
  assign io_wt_actv_data_0_0 = wt_actv_data_out_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_1 = wt_actv_data_out_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_2 = wt_actv_data_out_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_3 = wt_actv_data_out_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_4 = wt_actv_data_out_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_5 = wt_actv_data_out_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_6 = wt_actv_data_out_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_7 = wt_actv_data_out_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_8 = wt_actv_data_out_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_9 = wt_actv_data_out_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_10 = wt_actv_data_out_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_11 = wt_actv_data_out_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_12 = wt_actv_data_out_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_13 = wt_actv_data_out_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_14 = wt_actv_data_out_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_15 = wt_actv_data_out_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_16 = wt_actv_data_out_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_17 = wt_actv_data_out_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_18 = wt_actv_data_out_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_19 = wt_actv_data_out_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_20 = wt_actv_data_out_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_21 = wt_actv_data_out_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_22 = wt_actv_data_out_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_23 = wt_actv_data_out_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_24 = wt_actv_data_out_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_25 = wt_actv_data_out_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_26 = wt_actv_data_out_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_27 = wt_actv_data_out_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_28 = wt_actv_data_out_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_29 = wt_actv_data_out_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_30 = wt_actv_data_out_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_31 = wt_actv_data_out_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_32 = wt_actv_data_out_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_33 = wt_actv_data_out_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_34 = wt_actv_data_out_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_35 = wt_actv_data_out_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_36 = wt_actv_data_out_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_37 = wt_actv_data_out_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_38 = wt_actv_data_out_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_39 = wt_actv_data_out_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_40 = wt_actv_data_out_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_41 = wt_actv_data_out_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_42 = wt_actv_data_out_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_43 = wt_actv_data_out_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_44 = wt_actv_data_out_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_45 = wt_actv_data_out_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_46 = wt_actv_data_out_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_47 = wt_actv_data_out_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_48 = wt_actv_data_out_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_49 = wt_actv_data_out_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_50 = wt_actv_data_out_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_51 = wt_actv_data_out_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_52 = wt_actv_data_out_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_53 = wt_actv_data_out_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_54 = wt_actv_data_out_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_55 = wt_actv_data_out_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_56 = wt_actv_data_out_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_57 = wt_actv_data_out_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_58 = wt_actv_data_out_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_59 = wt_actv_data_out_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_60 = wt_actv_data_out_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_61 = wt_actv_data_out_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_62 = wt_actv_data_out_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_63 = wt_actv_data_out_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_64 = wt_actv_data_out_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_65 = wt_actv_data_out_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_66 = wt_actv_data_out_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_67 = wt_actv_data_out_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_68 = wt_actv_data_out_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_69 = wt_actv_data_out_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_70 = wt_actv_data_out_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_71 = wt_actv_data_out_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_72 = wt_actv_data_out_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_73 = wt_actv_data_out_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_74 = wt_actv_data_out_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_75 = wt_actv_data_out_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_76 = wt_actv_data_out_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_77 = wt_actv_data_out_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_78 = wt_actv_data_out_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_79 = wt_actv_data_out_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_80 = wt_actv_data_out_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_81 = wt_actv_data_out_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_82 = wt_actv_data_out_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_83 = wt_actv_data_out_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_84 = wt_actv_data_out_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_85 = wt_actv_data_out_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_86 = wt_actv_data_out_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_87 = wt_actv_data_out_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_88 = wt_actv_data_out_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_89 = wt_actv_data_out_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_90 = wt_actv_data_out_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_91 = wt_actv_data_out_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_92 = wt_actv_data_out_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_93 = wt_actv_data_out_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_94 = wt_actv_data_out_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_95 = wt_actv_data_out_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_96 = wt_actv_data_out_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_97 = wt_actv_data_out_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_98 = wt_actv_data_out_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_99 = wt_actv_data_out_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_100 = wt_actv_data_out_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_101 = wt_actv_data_out_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_102 = wt_actv_data_out_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_103 = wt_actv_data_out_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_104 = wt_actv_data_out_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_105 = wt_actv_data_out_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_106 = wt_actv_data_out_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_107 = wt_actv_data_out_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_108 = wt_actv_data_out_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_109 = wt_actv_data_out_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_110 = wt_actv_data_out_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_111 = wt_actv_data_out_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_112 = wt_actv_data_out_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_113 = wt_actv_data_out_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_114 = wt_actv_data_out_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_115 = wt_actv_data_out_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_116 = wt_actv_data_out_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_117 = wt_actv_data_out_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_118 = wt_actv_data_out_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_119 = wt_actv_data_out_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_120 = wt_actv_data_out_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_121 = wt_actv_data_out_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_122 = wt_actv_data_out_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_123 = wt_actv_data_out_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_124 = wt_actv_data_out_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_125 = wt_actv_data_out_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_126 = wt_actv_data_out_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_data_0_127 = wt_actv_data_out_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 183:21]
  assign io_wt_actv_nz_0_0 = wt_actv_nz_out_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_1 = wt_actv_nz_out_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_2 = wt_actv_nz_out_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_3 = wt_actv_nz_out_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_4 = wt_actv_nz_out_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_5 = wt_actv_nz_out_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_6 = wt_actv_nz_out_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_7 = wt_actv_nz_out_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_8 = wt_actv_nz_out_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_9 = wt_actv_nz_out_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_10 = wt_actv_nz_out_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_11 = wt_actv_nz_out_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_12 = wt_actv_nz_out_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_13 = wt_actv_nz_out_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_14 = wt_actv_nz_out_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_15 = wt_actv_nz_out_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_16 = wt_actv_nz_out_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_17 = wt_actv_nz_out_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_18 = wt_actv_nz_out_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_19 = wt_actv_nz_out_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_20 = wt_actv_nz_out_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_21 = wt_actv_nz_out_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_22 = wt_actv_nz_out_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_23 = wt_actv_nz_out_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_24 = wt_actv_nz_out_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_25 = wt_actv_nz_out_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_26 = wt_actv_nz_out_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_27 = wt_actv_nz_out_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_28 = wt_actv_nz_out_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_29 = wt_actv_nz_out_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_30 = wt_actv_nz_out_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_31 = wt_actv_nz_out_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_32 = wt_actv_nz_out_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_33 = wt_actv_nz_out_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_34 = wt_actv_nz_out_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_35 = wt_actv_nz_out_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_36 = wt_actv_nz_out_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_37 = wt_actv_nz_out_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_38 = wt_actv_nz_out_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_39 = wt_actv_nz_out_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_40 = wt_actv_nz_out_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_41 = wt_actv_nz_out_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_42 = wt_actv_nz_out_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_43 = wt_actv_nz_out_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_44 = wt_actv_nz_out_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_45 = wt_actv_nz_out_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_46 = wt_actv_nz_out_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_47 = wt_actv_nz_out_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_48 = wt_actv_nz_out_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_49 = wt_actv_nz_out_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_50 = wt_actv_nz_out_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_51 = wt_actv_nz_out_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_52 = wt_actv_nz_out_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_53 = wt_actv_nz_out_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_54 = wt_actv_nz_out_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_55 = wt_actv_nz_out_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_56 = wt_actv_nz_out_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_57 = wt_actv_nz_out_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_58 = wt_actv_nz_out_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_59 = wt_actv_nz_out_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_60 = wt_actv_nz_out_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_61 = wt_actv_nz_out_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_62 = wt_actv_nz_out_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_63 = wt_actv_nz_out_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_64 = wt_actv_nz_out_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_65 = wt_actv_nz_out_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_66 = wt_actv_nz_out_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_67 = wt_actv_nz_out_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_68 = wt_actv_nz_out_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_69 = wt_actv_nz_out_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_70 = wt_actv_nz_out_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_71 = wt_actv_nz_out_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_72 = wt_actv_nz_out_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_73 = wt_actv_nz_out_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_74 = wt_actv_nz_out_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_75 = wt_actv_nz_out_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_76 = wt_actv_nz_out_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_77 = wt_actv_nz_out_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_78 = wt_actv_nz_out_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_79 = wt_actv_nz_out_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_80 = wt_actv_nz_out_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_81 = wt_actv_nz_out_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_82 = wt_actv_nz_out_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_83 = wt_actv_nz_out_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_84 = wt_actv_nz_out_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_85 = wt_actv_nz_out_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_86 = wt_actv_nz_out_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_87 = wt_actv_nz_out_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_88 = wt_actv_nz_out_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_89 = wt_actv_nz_out_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_90 = wt_actv_nz_out_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_91 = wt_actv_nz_out_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_92 = wt_actv_nz_out_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_93 = wt_actv_nz_out_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_94 = wt_actv_nz_out_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_95 = wt_actv_nz_out_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_96 = wt_actv_nz_out_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_97 = wt_actv_nz_out_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_98 = wt_actv_nz_out_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_99 = wt_actv_nz_out_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_100 = wt_actv_nz_out_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_101 = wt_actv_nz_out_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_102 = wt_actv_nz_out_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_103 = wt_actv_nz_out_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_104 = wt_actv_nz_out_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_105 = wt_actv_nz_out_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_106 = wt_actv_nz_out_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_107 = wt_actv_nz_out_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_108 = wt_actv_nz_out_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_109 = wt_actv_nz_out_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_110 = wt_actv_nz_out_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_111 = wt_actv_nz_out_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_112 = wt_actv_nz_out_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_113 = wt_actv_nz_out_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_114 = wt_actv_nz_out_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_115 = wt_actv_nz_out_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_116 = wt_actv_nz_out_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_117 = wt_actv_nz_out_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_118 = wt_actv_nz_out_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_119 = wt_actv_nz_out_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_120 = wt_actv_nz_out_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_121 = wt_actv_nz_out_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_122 = wt_actv_nz_out_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_123 = wt_actv_nz_out_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_124 = wt_actv_nz_out_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_125 = wt_actv_nz_out_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_126 = wt_actv_nz_out_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_nz_0_127 = wt_actv_nz_out_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 184:19]
  assign io_wt_actv_pvld_0_0 = wt_actv_pvld_out_0_0; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_1 = wt_actv_pvld_out_0_1; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_2 = wt_actv_pvld_out_0_2; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_3 = wt_actv_pvld_out_0_3; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_4 = wt_actv_pvld_out_0_4; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_5 = wt_actv_pvld_out_0_5; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_6 = wt_actv_pvld_out_0_6; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_7 = wt_actv_pvld_out_0_7; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_8 = wt_actv_pvld_out_0_8; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_9 = wt_actv_pvld_out_0_9; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_10 = wt_actv_pvld_out_0_10; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_11 = wt_actv_pvld_out_0_11; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_12 = wt_actv_pvld_out_0_12; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_13 = wt_actv_pvld_out_0_13; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_14 = wt_actv_pvld_out_0_14; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_15 = wt_actv_pvld_out_0_15; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_16 = wt_actv_pvld_out_0_16; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_17 = wt_actv_pvld_out_0_17; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_18 = wt_actv_pvld_out_0_18; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_19 = wt_actv_pvld_out_0_19; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_20 = wt_actv_pvld_out_0_20; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_21 = wt_actv_pvld_out_0_21; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_22 = wt_actv_pvld_out_0_22; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_23 = wt_actv_pvld_out_0_23; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_24 = wt_actv_pvld_out_0_24; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_25 = wt_actv_pvld_out_0_25; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_26 = wt_actv_pvld_out_0_26; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_27 = wt_actv_pvld_out_0_27; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_28 = wt_actv_pvld_out_0_28; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_29 = wt_actv_pvld_out_0_29; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_30 = wt_actv_pvld_out_0_30; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_31 = wt_actv_pvld_out_0_31; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_32 = wt_actv_pvld_out_0_32; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_33 = wt_actv_pvld_out_0_33; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_34 = wt_actv_pvld_out_0_34; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_35 = wt_actv_pvld_out_0_35; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_36 = wt_actv_pvld_out_0_36; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_37 = wt_actv_pvld_out_0_37; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_38 = wt_actv_pvld_out_0_38; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_39 = wt_actv_pvld_out_0_39; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_40 = wt_actv_pvld_out_0_40; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_41 = wt_actv_pvld_out_0_41; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_42 = wt_actv_pvld_out_0_42; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_43 = wt_actv_pvld_out_0_43; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_44 = wt_actv_pvld_out_0_44; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_45 = wt_actv_pvld_out_0_45; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_46 = wt_actv_pvld_out_0_46; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_47 = wt_actv_pvld_out_0_47; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_48 = wt_actv_pvld_out_0_48; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_49 = wt_actv_pvld_out_0_49; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_50 = wt_actv_pvld_out_0_50; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_51 = wt_actv_pvld_out_0_51; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_52 = wt_actv_pvld_out_0_52; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_53 = wt_actv_pvld_out_0_53; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_54 = wt_actv_pvld_out_0_54; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_55 = wt_actv_pvld_out_0_55; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_56 = wt_actv_pvld_out_0_56; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_57 = wt_actv_pvld_out_0_57; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_58 = wt_actv_pvld_out_0_58; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_59 = wt_actv_pvld_out_0_59; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_60 = wt_actv_pvld_out_0_60; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_61 = wt_actv_pvld_out_0_61; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_62 = wt_actv_pvld_out_0_62; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_63 = wt_actv_pvld_out_0_63; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_64 = wt_actv_pvld_out_0_64; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_65 = wt_actv_pvld_out_0_65; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_66 = wt_actv_pvld_out_0_66; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_67 = wt_actv_pvld_out_0_67; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_68 = wt_actv_pvld_out_0_68; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_69 = wt_actv_pvld_out_0_69; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_70 = wt_actv_pvld_out_0_70; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_71 = wt_actv_pvld_out_0_71; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_72 = wt_actv_pvld_out_0_72; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_73 = wt_actv_pvld_out_0_73; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_74 = wt_actv_pvld_out_0_74; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_75 = wt_actv_pvld_out_0_75; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_76 = wt_actv_pvld_out_0_76; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_77 = wt_actv_pvld_out_0_77; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_78 = wt_actv_pvld_out_0_78; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_79 = wt_actv_pvld_out_0_79; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_80 = wt_actv_pvld_out_0_80; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_81 = wt_actv_pvld_out_0_81; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_82 = wt_actv_pvld_out_0_82; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_83 = wt_actv_pvld_out_0_83; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_84 = wt_actv_pvld_out_0_84; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_85 = wt_actv_pvld_out_0_85; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_86 = wt_actv_pvld_out_0_86; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_87 = wt_actv_pvld_out_0_87; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_88 = wt_actv_pvld_out_0_88; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_89 = wt_actv_pvld_out_0_89; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_90 = wt_actv_pvld_out_0_90; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_91 = wt_actv_pvld_out_0_91; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_92 = wt_actv_pvld_out_0_92; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_93 = wt_actv_pvld_out_0_93; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_94 = wt_actv_pvld_out_0_94; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_95 = wt_actv_pvld_out_0_95; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_96 = wt_actv_pvld_out_0_96; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_97 = wt_actv_pvld_out_0_97; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_98 = wt_actv_pvld_out_0_98; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_99 = wt_actv_pvld_out_0_99; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_100 = wt_actv_pvld_out_0_100; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_101 = wt_actv_pvld_out_0_101; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_102 = wt_actv_pvld_out_0_102; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_103 = wt_actv_pvld_out_0_103; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_104 = wt_actv_pvld_out_0_104; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_105 = wt_actv_pvld_out_0_105; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_106 = wt_actv_pvld_out_0_106; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_107 = wt_actv_pvld_out_0_107; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_108 = wt_actv_pvld_out_0_108; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_109 = wt_actv_pvld_out_0_109; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_110 = wt_actv_pvld_out_0_110; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_111 = wt_actv_pvld_out_0_111; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_112 = wt_actv_pvld_out_0_112; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_113 = wt_actv_pvld_out_0_113; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_114 = wt_actv_pvld_out_0_114; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_115 = wt_actv_pvld_out_0_115; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_116 = wt_actv_pvld_out_0_116; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_117 = wt_actv_pvld_out_0_117; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_118 = wt_actv_pvld_out_0_118; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_119 = wt_actv_pvld_out_0_119; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_120 = wt_actv_pvld_out_0_120; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_121 = wt_actv_pvld_out_0_121; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_122 = wt_actv_pvld_out_0_122; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_123 = wt_actv_pvld_out_0_123; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_124 = wt_actv_pvld_out_0_124; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_125 = wt_actv_pvld_out_0_125; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_126 = wt_actv_pvld_out_0_126; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
  assign io_wt_actv_pvld_0_127 = wt_actv_pvld_out_0_127; // @[NV_NVDLA_CMAC_CORE_active.scala 182:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wt_pre_nz_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  wt_pre_nz_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  wt_pre_nz_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  wt_pre_nz_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  wt_pre_nz_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  wt_pre_nz_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  wt_pre_nz_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  wt_pre_nz_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wt_pre_nz_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wt_pre_nz_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wt_pre_nz_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wt_pre_nz_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wt_pre_nz_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wt_pre_nz_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wt_pre_nz_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  wt_pre_nz_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  wt_pre_nz_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  wt_pre_nz_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wt_pre_nz_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  wt_pre_nz_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  wt_pre_nz_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  wt_pre_nz_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  wt_pre_nz_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  wt_pre_nz_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  wt_pre_nz_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  wt_pre_nz_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  wt_pre_nz_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  wt_pre_nz_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  wt_pre_nz_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  wt_pre_nz_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  wt_pre_nz_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  wt_pre_nz_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  wt_pre_nz_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wt_pre_nz_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  wt_pre_nz_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wt_pre_nz_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wt_pre_nz_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  wt_pre_nz_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  wt_pre_nz_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  wt_pre_nz_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  wt_pre_nz_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  wt_pre_nz_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  wt_pre_nz_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  wt_pre_nz_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  wt_pre_nz_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  wt_pre_nz_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  wt_pre_nz_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  wt_pre_nz_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  wt_pre_nz_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  wt_pre_nz_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  wt_pre_nz_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  wt_pre_nz_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  wt_pre_nz_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  wt_pre_nz_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  wt_pre_nz_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  wt_pre_nz_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  wt_pre_nz_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  wt_pre_nz_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  wt_pre_nz_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  wt_pre_nz_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  wt_pre_nz_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  wt_pre_nz_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  wt_pre_nz_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  wt_pre_nz_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  wt_pre_nz_64 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  wt_pre_nz_65 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  wt_pre_nz_66 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  wt_pre_nz_67 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  wt_pre_nz_68 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  wt_pre_nz_69 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  wt_pre_nz_70 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  wt_pre_nz_71 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  wt_pre_nz_72 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  wt_pre_nz_73 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  wt_pre_nz_74 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  wt_pre_nz_75 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  wt_pre_nz_76 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  wt_pre_nz_77 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  wt_pre_nz_78 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  wt_pre_nz_79 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  wt_pre_nz_80 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  wt_pre_nz_81 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  wt_pre_nz_82 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  wt_pre_nz_83 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  wt_pre_nz_84 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  wt_pre_nz_85 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  wt_pre_nz_86 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  wt_pre_nz_87 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  wt_pre_nz_88 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  wt_pre_nz_89 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  wt_pre_nz_90 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  wt_pre_nz_91 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  wt_pre_nz_92 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  wt_pre_nz_93 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  wt_pre_nz_94 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  wt_pre_nz_95 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  wt_pre_nz_96 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  wt_pre_nz_97 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  wt_pre_nz_98 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  wt_pre_nz_99 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  wt_pre_nz_100 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  wt_pre_nz_101 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  wt_pre_nz_102 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  wt_pre_nz_103 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  wt_pre_nz_104 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  wt_pre_nz_105 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  wt_pre_nz_106 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  wt_pre_nz_107 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  wt_pre_nz_108 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  wt_pre_nz_109 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  wt_pre_nz_110 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  wt_pre_nz_111 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  wt_pre_nz_112 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  wt_pre_nz_113 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  wt_pre_nz_114 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  wt_pre_nz_115 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  wt_pre_nz_116 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  wt_pre_nz_117 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  wt_pre_nz_118 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  wt_pre_nz_119 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  wt_pre_nz_120 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  wt_pre_nz_121 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  wt_pre_nz_122 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  wt_pre_nz_123 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  wt_pre_nz_124 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  wt_pre_nz_125 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  wt_pre_nz_126 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  wt_pre_nz_127 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  wt_pre_data_0 = _RAND_128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  wt_pre_data_1 = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  wt_pre_data_2 = _RAND_130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  wt_pre_data_3 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  wt_pre_data_4 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  wt_pre_data_5 = _RAND_133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  wt_pre_data_6 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  wt_pre_data_7 = _RAND_135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  wt_pre_data_8 = _RAND_136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  wt_pre_data_9 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  wt_pre_data_10 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  wt_pre_data_11 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  wt_pre_data_12 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  wt_pre_data_13 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  wt_pre_data_14 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  wt_pre_data_15 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  wt_pre_data_16 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  wt_pre_data_17 = _RAND_145[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  wt_pre_data_18 = _RAND_146[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  wt_pre_data_19 = _RAND_147[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  wt_pre_data_20 = _RAND_148[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  wt_pre_data_21 = _RAND_149[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  wt_pre_data_22 = _RAND_150[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  wt_pre_data_23 = _RAND_151[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  wt_pre_data_24 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  wt_pre_data_25 = _RAND_153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  wt_pre_data_26 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  wt_pre_data_27 = _RAND_155[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  wt_pre_data_28 = _RAND_156[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  wt_pre_data_29 = _RAND_157[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  wt_pre_data_30 = _RAND_158[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  wt_pre_data_31 = _RAND_159[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  wt_pre_data_32 = _RAND_160[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  wt_pre_data_33 = _RAND_161[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  wt_pre_data_34 = _RAND_162[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  wt_pre_data_35 = _RAND_163[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  wt_pre_data_36 = _RAND_164[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  wt_pre_data_37 = _RAND_165[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  wt_pre_data_38 = _RAND_166[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  wt_pre_data_39 = _RAND_167[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  wt_pre_data_40 = _RAND_168[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  wt_pre_data_41 = _RAND_169[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  wt_pre_data_42 = _RAND_170[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  wt_pre_data_43 = _RAND_171[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  wt_pre_data_44 = _RAND_172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  wt_pre_data_45 = _RAND_173[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  wt_pre_data_46 = _RAND_174[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  wt_pre_data_47 = _RAND_175[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  wt_pre_data_48 = _RAND_176[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  wt_pre_data_49 = _RAND_177[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  wt_pre_data_50 = _RAND_178[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  wt_pre_data_51 = _RAND_179[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  wt_pre_data_52 = _RAND_180[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  wt_pre_data_53 = _RAND_181[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  wt_pre_data_54 = _RAND_182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  wt_pre_data_55 = _RAND_183[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  wt_pre_data_56 = _RAND_184[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  wt_pre_data_57 = _RAND_185[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  wt_pre_data_58 = _RAND_186[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  wt_pre_data_59 = _RAND_187[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  wt_pre_data_60 = _RAND_188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  wt_pre_data_61 = _RAND_189[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  wt_pre_data_62 = _RAND_190[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  wt_pre_data_63 = _RAND_191[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  wt_pre_data_64 = _RAND_192[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  wt_pre_data_65 = _RAND_193[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  wt_pre_data_66 = _RAND_194[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  wt_pre_data_67 = _RAND_195[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  wt_pre_data_68 = _RAND_196[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  wt_pre_data_69 = _RAND_197[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  wt_pre_data_70 = _RAND_198[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  wt_pre_data_71 = _RAND_199[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  wt_pre_data_72 = _RAND_200[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  wt_pre_data_73 = _RAND_201[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  wt_pre_data_74 = _RAND_202[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  wt_pre_data_75 = _RAND_203[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  wt_pre_data_76 = _RAND_204[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  wt_pre_data_77 = _RAND_205[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  wt_pre_data_78 = _RAND_206[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  wt_pre_data_79 = _RAND_207[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  wt_pre_data_80 = _RAND_208[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  wt_pre_data_81 = _RAND_209[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  wt_pre_data_82 = _RAND_210[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  wt_pre_data_83 = _RAND_211[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  wt_pre_data_84 = _RAND_212[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  wt_pre_data_85 = _RAND_213[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  wt_pre_data_86 = _RAND_214[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  wt_pre_data_87 = _RAND_215[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  wt_pre_data_88 = _RAND_216[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  wt_pre_data_89 = _RAND_217[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  wt_pre_data_90 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  wt_pre_data_91 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  wt_pre_data_92 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  wt_pre_data_93 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  wt_pre_data_94 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  wt_pre_data_95 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  wt_pre_data_96 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  wt_pre_data_97 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  wt_pre_data_98 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  wt_pre_data_99 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  wt_pre_data_100 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  wt_pre_data_101 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  wt_pre_data_102 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  wt_pre_data_103 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  wt_pre_data_104 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  wt_pre_data_105 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  wt_pre_data_106 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  wt_pre_data_107 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  wt_pre_data_108 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  wt_pre_data_109 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  wt_pre_data_110 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  wt_pre_data_111 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  wt_pre_data_112 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  wt_pre_data_113 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  wt_pre_data_114 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  wt_pre_data_115 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  wt_pre_data_116 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  wt_pre_data_117 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  wt_pre_data_118 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  wt_pre_data_119 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  wt_pre_data_120 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  wt_pre_data_121 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  wt_pre_data_122 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  wt_pre_data_123 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  wt_pre_data_124 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  wt_pre_data_125 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  wt_pre_data_126 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  wt_pre_data_127 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  wt_pre_sel_0 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  dat_pre_nz_0 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  dat_pre_nz_1 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  dat_pre_nz_2 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  dat_pre_nz_3 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  dat_pre_nz_4 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  dat_pre_nz_5 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  dat_pre_nz_6 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  dat_pre_nz_7 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  dat_pre_nz_8 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  dat_pre_nz_9 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  dat_pre_nz_10 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  dat_pre_nz_11 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  dat_pre_nz_12 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  dat_pre_nz_13 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  dat_pre_nz_14 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  dat_pre_nz_15 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  dat_pre_nz_16 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  dat_pre_nz_17 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  dat_pre_nz_18 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  dat_pre_nz_19 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  dat_pre_nz_20 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  dat_pre_nz_21 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  dat_pre_nz_22 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  dat_pre_nz_23 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  dat_pre_nz_24 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  dat_pre_nz_25 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  dat_pre_nz_26 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  dat_pre_nz_27 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  dat_pre_nz_28 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  dat_pre_nz_29 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  dat_pre_nz_30 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  dat_pre_nz_31 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  dat_pre_nz_32 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  dat_pre_nz_33 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  dat_pre_nz_34 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  dat_pre_nz_35 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  dat_pre_nz_36 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  dat_pre_nz_37 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  dat_pre_nz_38 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  dat_pre_nz_39 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  dat_pre_nz_40 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  dat_pre_nz_41 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  dat_pre_nz_42 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  dat_pre_nz_43 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  dat_pre_nz_44 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  dat_pre_nz_45 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  dat_pre_nz_46 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  dat_pre_nz_47 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  dat_pre_nz_48 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  dat_pre_nz_49 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  dat_pre_nz_50 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  dat_pre_nz_51 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  dat_pre_nz_52 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  dat_pre_nz_53 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  dat_pre_nz_54 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  dat_pre_nz_55 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  dat_pre_nz_56 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  dat_pre_nz_57 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  dat_pre_nz_58 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  dat_pre_nz_59 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  dat_pre_nz_60 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  dat_pre_nz_61 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  dat_pre_nz_62 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  dat_pre_nz_63 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  dat_pre_nz_64 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  dat_pre_nz_65 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  dat_pre_nz_66 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  dat_pre_nz_67 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  dat_pre_nz_68 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  dat_pre_nz_69 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  dat_pre_nz_70 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  dat_pre_nz_71 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  dat_pre_nz_72 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  dat_pre_nz_73 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  dat_pre_nz_74 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  dat_pre_nz_75 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  dat_pre_nz_76 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  dat_pre_nz_77 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  dat_pre_nz_78 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  dat_pre_nz_79 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  dat_pre_nz_80 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  dat_pre_nz_81 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  dat_pre_nz_82 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  dat_pre_nz_83 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  dat_pre_nz_84 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  dat_pre_nz_85 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  dat_pre_nz_86 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  dat_pre_nz_87 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  dat_pre_nz_88 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  dat_pre_nz_89 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  dat_pre_nz_90 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  dat_pre_nz_91 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  dat_pre_nz_92 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  dat_pre_nz_93 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  dat_pre_nz_94 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  dat_pre_nz_95 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  dat_pre_nz_96 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  dat_pre_nz_97 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  dat_pre_nz_98 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  dat_pre_nz_99 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  dat_pre_nz_100 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  dat_pre_nz_101 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  dat_pre_nz_102 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  dat_pre_nz_103 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  dat_pre_nz_104 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  dat_pre_nz_105 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  dat_pre_nz_106 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  dat_pre_nz_107 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  dat_pre_nz_108 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  dat_pre_nz_109 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  dat_pre_nz_110 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  dat_pre_nz_111 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  dat_pre_nz_112 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  dat_pre_nz_113 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  dat_pre_nz_114 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  dat_pre_nz_115 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  dat_pre_nz_116 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  dat_pre_nz_117 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  dat_pre_nz_118 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  dat_pre_nz_119 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  dat_pre_nz_120 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  dat_pre_nz_121 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  dat_pre_nz_122 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  dat_pre_nz_123 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  dat_pre_nz_124 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  dat_pre_nz_125 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  dat_pre_nz_126 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  dat_pre_nz_127 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  dat_pre_data_0 = _RAND_385[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  dat_pre_data_1 = _RAND_386[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  dat_pre_data_2 = _RAND_387[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  dat_pre_data_3 = _RAND_388[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  dat_pre_data_4 = _RAND_389[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  dat_pre_data_5 = _RAND_390[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  dat_pre_data_6 = _RAND_391[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  dat_pre_data_7 = _RAND_392[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  dat_pre_data_8 = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  dat_pre_data_9 = _RAND_394[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  dat_pre_data_10 = _RAND_395[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  dat_pre_data_11 = _RAND_396[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  dat_pre_data_12 = _RAND_397[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  dat_pre_data_13 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  dat_pre_data_14 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  dat_pre_data_15 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  dat_pre_data_16 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  dat_pre_data_17 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  dat_pre_data_18 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  dat_pre_data_19 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  dat_pre_data_20 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  dat_pre_data_21 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  dat_pre_data_22 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  dat_pre_data_23 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  dat_pre_data_24 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  dat_pre_data_25 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  dat_pre_data_26 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  dat_pre_data_27 = _RAND_412[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  dat_pre_data_28 = _RAND_413[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  dat_pre_data_29 = _RAND_414[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  dat_pre_data_30 = _RAND_415[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  dat_pre_data_31 = _RAND_416[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  dat_pre_data_32 = _RAND_417[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  dat_pre_data_33 = _RAND_418[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  dat_pre_data_34 = _RAND_419[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  dat_pre_data_35 = _RAND_420[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  dat_pre_data_36 = _RAND_421[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  dat_pre_data_37 = _RAND_422[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  dat_pre_data_38 = _RAND_423[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  dat_pre_data_39 = _RAND_424[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  dat_pre_data_40 = _RAND_425[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  dat_pre_data_41 = _RAND_426[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  dat_pre_data_42 = _RAND_427[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  dat_pre_data_43 = _RAND_428[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  dat_pre_data_44 = _RAND_429[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  dat_pre_data_45 = _RAND_430[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  dat_pre_data_46 = _RAND_431[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  dat_pre_data_47 = _RAND_432[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  dat_pre_data_48 = _RAND_433[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  dat_pre_data_49 = _RAND_434[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  dat_pre_data_50 = _RAND_435[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  dat_pre_data_51 = _RAND_436[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  dat_pre_data_52 = _RAND_437[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  dat_pre_data_53 = _RAND_438[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  dat_pre_data_54 = _RAND_439[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  dat_pre_data_55 = _RAND_440[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  dat_pre_data_56 = _RAND_441[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  dat_pre_data_57 = _RAND_442[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  dat_pre_data_58 = _RAND_443[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  dat_pre_data_59 = _RAND_444[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  dat_pre_data_60 = _RAND_445[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  dat_pre_data_61 = _RAND_446[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  dat_pre_data_62 = _RAND_447[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  dat_pre_data_63 = _RAND_448[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  dat_pre_data_64 = _RAND_449[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  dat_pre_data_65 = _RAND_450[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  dat_pre_data_66 = _RAND_451[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  dat_pre_data_67 = _RAND_452[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  dat_pre_data_68 = _RAND_453[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  dat_pre_data_69 = _RAND_454[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  dat_pre_data_70 = _RAND_455[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  dat_pre_data_71 = _RAND_456[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  dat_pre_data_72 = _RAND_457[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  dat_pre_data_73 = _RAND_458[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  dat_pre_data_74 = _RAND_459[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  dat_pre_data_75 = _RAND_460[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  dat_pre_data_76 = _RAND_461[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  dat_pre_data_77 = _RAND_462[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  dat_pre_data_78 = _RAND_463[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  dat_pre_data_79 = _RAND_464[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  dat_pre_data_80 = _RAND_465[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  dat_pre_data_81 = _RAND_466[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  dat_pre_data_82 = _RAND_467[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  dat_pre_data_83 = _RAND_468[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  dat_pre_data_84 = _RAND_469[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  dat_pre_data_85 = _RAND_470[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  dat_pre_data_86 = _RAND_471[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  dat_pre_data_87 = _RAND_472[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  dat_pre_data_88 = _RAND_473[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  dat_pre_data_89 = _RAND_474[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  dat_pre_data_90 = _RAND_475[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  dat_pre_data_91 = _RAND_476[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  dat_pre_data_92 = _RAND_477[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  dat_pre_data_93 = _RAND_478[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  dat_pre_data_94 = _RAND_479[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  dat_pre_data_95 = _RAND_480[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  dat_pre_data_96 = _RAND_481[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  dat_pre_data_97 = _RAND_482[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  dat_pre_data_98 = _RAND_483[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  dat_pre_data_99 = _RAND_484[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  dat_pre_data_100 = _RAND_485[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  dat_pre_data_101 = _RAND_486[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  dat_pre_data_102 = _RAND_487[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  dat_pre_data_103 = _RAND_488[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  dat_pre_data_104 = _RAND_489[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  dat_pre_data_105 = _RAND_490[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  dat_pre_data_106 = _RAND_491[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  dat_pre_data_107 = _RAND_492[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  dat_pre_data_108 = _RAND_493[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  dat_pre_data_109 = _RAND_494[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  dat_pre_data_110 = _RAND_495[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  dat_pre_data_111 = _RAND_496[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  dat_pre_data_112 = _RAND_497[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  dat_pre_data_113 = _RAND_498[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  dat_pre_data_114 = _RAND_499[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  dat_pre_data_115 = _RAND_500[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  dat_pre_data_116 = _RAND_501[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  dat_pre_data_117 = _RAND_502[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  dat_pre_data_118 = _RAND_503[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  dat_pre_data_119 = _RAND_504[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  dat_pre_data_120 = _RAND_505[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  dat_pre_data_121 = _RAND_506[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  dat_pre_data_122 = _RAND_507[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  dat_pre_data_123 = _RAND_508[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  dat_pre_data_124 = _RAND_509[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  dat_pre_data_125 = _RAND_510[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  dat_pre_data_126 = _RAND_511[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  dat_pre_data_127 = _RAND_512[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  dat_pre_pvld = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  dat_pre_stripe_st_out_0 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  dat_pre_stripe_end_out_0 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  wt_sd_pvld_0 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  wt_sd_nz_0_0 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  wt_sd_nz_0_1 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  wt_sd_nz_0_2 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  wt_sd_nz_0_3 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  wt_sd_nz_0_4 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  wt_sd_nz_0_5 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  wt_sd_nz_0_6 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  wt_sd_nz_0_7 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  wt_sd_nz_0_8 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  wt_sd_nz_0_9 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  wt_sd_nz_0_10 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  wt_sd_nz_0_11 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  wt_sd_nz_0_12 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  wt_sd_nz_0_13 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  wt_sd_nz_0_14 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  wt_sd_nz_0_15 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  wt_sd_nz_0_16 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  wt_sd_nz_0_17 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  wt_sd_nz_0_18 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  wt_sd_nz_0_19 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  wt_sd_nz_0_20 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  wt_sd_nz_0_21 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  wt_sd_nz_0_22 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  wt_sd_nz_0_23 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  wt_sd_nz_0_24 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  wt_sd_nz_0_25 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  wt_sd_nz_0_26 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  wt_sd_nz_0_27 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  wt_sd_nz_0_28 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  wt_sd_nz_0_29 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  wt_sd_nz_0_30 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  wt_sd_nz_0_31 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  wt_sd_nz_0_32 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  wt_sd_nz_0_33 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  wt_sd_nz_0_34 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  wt_sd_nz_0_35 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  wt_sd_nz_0_36 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  wt_sd_nz_0_37 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  wt_sd_nz_0_38 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  wt_sd_nz_0_39 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  wt_sd_nz_0_40 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  wt_sd_nz_0_41 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  wt_sd_nz_0_42 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  wt_sd_nz_0_43 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  wt_sd_nz_0_44 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  wt_sd_nz_0_45 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  wt_sd_nz_0_46 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  wt_sd_nz_0_47 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  wt_sd_nz_0_48 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  wt_sd_nz_0_49 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  wt_sd_nz_0_50 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  wt_sd_nz_0_51 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  wt_sd_nz_0_52 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  wt_sd_nz_0_53 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  wt_sd_nz_0_54 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  wt_sd_nz_0_55 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  wt_sd_nz_0_56 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  wt_sd_nz_0_57 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  wt_sd_nz_0_58 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  wt_sd_nz_0_59 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  wt_sd_nz_0_60 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  wt_sd_nz_0_61 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  wt_sd_nz_0_62 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  wt_sd_nz_0_63 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  wt_sd_nz_0_64 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  wt_sd_nz_0_65 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  wt_sd_nz_0_66 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  wt_sd_nz_0_67 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  wt_sd_nz_0_68 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  wt_sd_nz_0_69 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  wt_sd_nz_0_70 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  wt_sd_nz_0_71 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  wt_sd_nz_0_72 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  wt_sd_nz_0_73 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  wt_sd_nz_0_74 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  wt_sd_nz_0_75 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  wt_sd_nz_0_76 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  wt_sd_nz_0_77 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  wt_sd_nz_0_78 = _RAND_595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  wt_sd_nz_0_79 = _RAND_596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  wt_sd_nz_0_80 = _RAND_597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  wt_sd_nz_0_81 = _RAND_598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  wt_sd_nz_0_82 = _RAND_599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  wt_sd_nz_0_83 = _RAND_600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  wt_sd_nz_0_84 = _RAND_601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  wt_sd_nz_0_85 = _RAND_602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  wt_sd_nz_0_86 = _RAND_603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  wt_sd_nz_0_87 = _RAND_604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  wt_sd_nz_0_88 = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  wt_sd_nz_0_89 = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  wt_sd_nz_0_90 = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  wt_sd_nz_0_91 = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  wt_sd_nz_0_92 = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  wt_sd_nz_0_93 = _RAND_610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  wt_sd_nz_0_94 = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  wt_sd_nz_0_95 = _RAND_612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  wt_sd_nz_0_96 = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  wt_sd_nz_0_97 = _RAND_614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  wt_sd_nz_0_98 = _RAND_615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  wt_sd_nz_0_99 = _RAND_616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  wt_sd_nz_0_100 = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  wt_sd_nz_0_101 = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  wt_sd_nz_0_102 = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  wt_sd_nz_0_103 = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  wt_sd_nz_0_104 = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  wt_sd_nz_0_105 = _RAND_622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  wt_sd_nz_0_106 = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  wt_sd_nz_0_107 = _RAND_624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  wt_sd_nz_0_108 = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  wt_sd_nz_0_109 = _RAND_626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  wt_sd_nz_0_110 = _RAND_627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  wt_sd_nz_0_111 = _RAND_628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  wt_sd_nz_0_112 = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  wt_sd_nz_0_113 = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  wt_sd_nz_0_114 = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  wt_sd_nz_0_115 = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  wt_sd_nz_0_116 = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  wt_sd_nz_0_117 = _RAND_634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  wt_sd_nz_0_118 = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  wt_sd_nz_0_119 = _RAND_636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  wt_sd_nz_0_120 = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  wt_sd_nz_0_121 = _RAND_638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  wt_sd_nz_0_122 = _RAND_639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  wt_sd_nz_0_123 = _RAND_640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  wt_sd_nz_0_124 = _RAND_641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  wt_sd_nz_0_125 = _RAND_642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  wt_sd_nz_0_126 = _RAND_643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  wt_sd_nz_0_127 = _RAND_644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  wt_sd_data_0_0 = _RAND_645[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  wt_sd_data_0_1 = _RAND_646[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  wt_sd_data_0_2 = _RAND_647[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  wt_sd_data_0_3 = _RAND_648[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  wt_sd_data_0_4 = _RAND_649[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  wt_sd_data_0_5 = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  wt_sd_data_0_6 = _RAND_651[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  wt_sd_data_0_7 = _RAND_652[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  wt_sd_data_0_8 = _RAND_653[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  wt_sd_data_0_9 = _RAND_654[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  wt_sd_data_0_10 = _RAND_655[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  wt_sd_data_0_11 = _RAND_656[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  wt_sd_data_0_12 = _RAND_657[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  wt_sd_data_0_13 = _RAND_658[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  wt_sd_data_0_14 = _RAND_659[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  wt_sd_data_0_15 = _RAND_660[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  wt_sd_data_0_16 = _RAND_661[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  wt_sd_data_0_17 = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  wt_sd_data_0_18 = _RAND_663[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  wt_sd_data_0_19 = _RAND_664[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  wt_sd_data_0_20 = _RAND_665[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  wt_sd_data_0_21 = _RAND_666[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  wt_sd_data_0_22 = _RAND_667[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  wt_sd_data_0_23 = _RAND_668[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  wt_sd_data_0_24 = _RAND_669[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  wt_sd_data_0_25 = _RAND_670[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  wt_sd_data_0_26 = _RAND_671[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  wt_sd_data_0_27 = _RAND_672[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  wt_sd_data_0_28 = _RAND_673[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  wt_sd_data_0_29 = _RAND_674[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  wt_sd_data_0_30 = _RAND_675[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  wt_sd_data_0_31 = _RAND_676[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  wt_sd_data_0_32 = _RAND_677[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  wt_sd_data_0_33 = _RAND_678[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  wt_sd_data_0_34 = _RAND_679[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  wt_sd_data_0_35 = _RAND_680[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  wt_sd_data_0_36 = _RAND_681[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  wt_sd_data_0_37 = _RAND_682[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  wt_sd_data_0_38 = _RAND_683[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  wt_sd_data_0_39 = _RAND_684[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  wt_sd_data_0_40 = _RAND_685[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  wt_sd_data_0_41 = _RAND_686[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  wt_sd_data_0_42 = _RAND_687[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  wt_sd_data_0_43 = _RAND_688[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  wt_sd_data_0_44 = _RAND_689[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  wt_sd_data_0_45 = _RAND_690[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  wt_sd_data_0_46 = _RAND_691[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  wt_sd_data_0_47 = _RAND_692[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  wt_sd_data_0_48 = _RAND_693[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  wt_sd_data_0_49 = _RAND_694[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  wt_sd_data_0_50 = _RAND_695[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  wt_sd_data_0_51 = _RAND_696[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  wt_sd_data_0_52 = _RAND_697[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  wt_sd_data_0_53 = _RAND_698[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  wt_sd_data_0_54 = _RAND_699[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  wt_sd_data_0_55 = _RAND_700[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  wt_sd_data_0_56 = _RAND_701[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  wt_sd_data_0_57 = _RAND_702[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  wt_sd_data_0_58 = _RAND_703[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  wt_sd_data_0_59 = _RAND_704[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  wt_sd_data_0_60 = _RAND_705[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  wt_sd_data_0_61 = _RAND_706[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  wt_sd_data_0_62 = _RAND_707[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  wt_sd_data_0_63 = _RAND_708[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  wt_sd_data_0_64 = _RAND_709[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  wt_sd_data_0_65 = _RAND_710[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  wt_sd_data_0_66 = _RAND_711[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  wt_sd_data_0_67 = _RAND_712[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  wt_sd_data_0_68 = _RAND_713[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  wt_sd_data_0_69 = _RAND_714[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  wt_sd_data_0_70 = _RAND_715[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  wt_sd_data_0_71 = _RAND_716[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  wt_sd_data_0_72 = _RAND_717[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  wt_sd_data_0_73 = _RAND_718[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  wt_sd_data_0_74 = _RAND_719[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  wt_sd_data_0_75 = _RAND_720[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  wt_sd_data_0_76 = _RAND_721[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  wt_sd_data_0_77 = _RAND_722[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  wt_sd_data_0_78 = _RAND_723[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  wt_sd_data_0_79 = _RAND_724[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  wt_sd_data_0_80 = _RAND_725[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  wt_sd_data_0_81 = _RAND_726[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  wt_sd_data_0_82 = _RAND_727[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  wt_sd_data_0_83 = _RAND_728[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  wt_sd_data_0_84 = _RAND_729[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  wt_sd_data_0_85 = _RAND_730[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  wt_sd_data_0_86 = _RAND_731[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  wt_sd_data_0_87 = _RAND_732[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  wt_sd_data_0_88 = _RAND_733[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  wt_sd_data_0_89 = _RAND_734[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  wt_sd_data_0_90 = _RAND_735[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  wt_sd_data_0_91 = _RAND_736[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  wt_sd_data_0_92 = _RAND_737[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  wt_sd_data_0_93 = _RAND_738[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  wt_sd_data_0_94 = _RAND_739[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  wt_sd_data_0_95 = _RAND_740[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  wt_sd_data_0_96 = _RAND_741[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  wt_sd_data_0_97 = _RAND_742[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  wt_sd_data_0_98 = _RAND_743[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  wt_sd_data_0_99 = _RAND_744[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  wt_sd_data_0_100 = _RAND_745[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  wt_sd_data_0_101 = _RAND_746[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  wt_sd_data_0_102 = _RAND_747[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  wt_sd_data_0_103 = _RAND_748[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  wt_sd_data_0_104 = _RAND_749[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  wt_sd_data_0_105 = _RAND_750[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  wt_sd_data_0_106 = _RAND_751[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  wt_sd_data_0_107 = _RAND_752[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  wt_sd_data_0_108 = _RAND_753[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  wt_sd_data_0_109 = _RAND_754[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  wt_sd_data_0_110 = _RAND_755[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  wt_sd_data_0_111 = _RAND_756[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  wt_sd_data_0_112 = _RAND_757[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  wt_sd_data_0_113 = _RAND_758[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  wt_sd_data_0_114 = _RAND_759[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  wt_sd_data_0_115 = _RAND_760[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  wt_sd_data_0_116 = _RAND_761[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  wt_sd_data_0_117 = _RAND_762[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  wt_sd_data_0_118 = _RAND_763[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  wt_sd_data_0_119 = _RAND_764[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  wt_sd_data_0_120 = _RAND_765[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  wt_sd_data_0_121 = _RAND_766[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  wt_sd_data_0_122 = _RAND_767[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  wt_sd_data_0_123 = _RAND_768[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  wt_sd_data_0_124 = _RAND_769[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  wt_sd_data_0_125 = _RAND_770[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  wt_sd_data_0_126 = _RAND_771[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  wt_sd_data_0_127 = _RAND_772[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  dat_actv_stripe_end_0 = _RAND_773[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  wt_actv_vld_0 = _RAND_774[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  wt_actv_pvld_out_0_0 = _RAND_775[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  wt_actv_pvld_out_0_1 = _RAND_776[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  wt_actv_pvld_out_0_2 = _RAND_777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  wt_actv_pvld_out_0_3 = _RAND_778[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  wt_actv_pvld_out_0_4 = _RAND_779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  wt_actv_pvld_out_0_5 = _RAND_780[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  wt_actv_pvld_out_0_6 = _RAND_781[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  wt_actv_pvld_out_0_7 = _RAND_782[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  wt_actv_pvld_out_0_8 = _RAND_783[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  wt_actv_pvld_out_0_9 = _RAND_784[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  wt_actv_pvld_out_0_10 = _RAND_785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  wt_actv_pvld_out_0_11 = _RAND_786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  wt_actv_pvld_out_0_12 = _RAND_787[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  wt_actv_pvld_out_0_13 = _RAND_788[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  wt_actv_pvld_out_0_14 = _RAND_789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  wt_actv_pvld_out_0_15 = _RAND_790[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  wt_actv_pvld_out_0_16 = _RAND_791[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  wt_actv_pvld_out_0_17 = _RAND_792[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  wt_actv_pvld_out_0_18 = _RAND_793[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  wt_actv_pvld_out_0_19 = _RAND_794[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  wt_actv_pvld_out_0_20 = _RAND_795[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  wt_actv_pvld_out_0_21 = _RAND_796[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  wt_actv_pvld_out_0_22 = _RAND_797[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  wt_actv_pvld_out_0_23 = _RAND_798[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  wt_actv_pvld_out_0_24 = _RAND_799[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  wt_actv_pvld_out_0_25 = _RAND_800[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  wt_actv_pvld_out_0_26 = _RAND_801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  wt_actv_pvld_out_0_27 = _RAND_802[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  wt_actv_pvld_out_0_28 = _RAND_803[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  wt_actv_pvld_out_0_29 = _RAND_804[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  wt_actv_pvld_out_0_30 = _RAND_805[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  wt_actv_pvld_out_0_31 = _RAND_806[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  wt_actv_pvld_out_0_32 = _RAND_807[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  wt_actv_pvld_out_0_33 = _RAND_808[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  wt_actv_pvld_out_0_34 = _RAND_809[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  wt_actv_pvld_out_0_35 = _RAND_810[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  wt_actv_pvld_out_0_36 = _RAND_811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  wt_actv_pvld_out_0_37 = _RAND_812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  wt_actv_pvld_out_0_38 = _RAND_813[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  wt_actv_pvld_out_0_39 = _RAND_814[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  wt_actv_pvld_out_0_40 = _RAND_815[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  wt_actv_pvld_out_0_41 = _RAND_816[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  wt_actv_pvld_out_0_42 = _RAND_817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  wt_actv_pvld_out_0_43 = _RAND_818[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  wt_actv_pvld_out_0_44 = _RAND_819[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  wt_actv_pvld_out_0_45 = _RAND_820[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  wt_actv_pvld_out_0_46 = _RAND_821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  wt_actv_pvld_out_0_47 = _RAND_822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  wt_actv_pvld_out_0_48 = _RAND_823[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  wt_actv_pvld_out_0_49 = _RAND_824[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  wt_actv_pvld_out_0_50 = _RAND_825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  wt_actv_pvld_out_0_51 = _RAND_826[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  wt_actv_pvld_out_0_52 = _RAND_827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  wt_actv_pvld_out_0_53 = _RAND_828[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  wt_actv_pvld_out_0_54 = _RAND_829[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  wt_actv_pvld_out_0_55 = _RAND_830[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  wt_actv_pvld_out_0_56 = _RAND_831[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  wt_actv_pvld_out_0_57 = _RAND_832[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  wt_actv_pvld_out_0_58 = _RAND_833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  wt_actv_pvld_out_0_59 = _RAND_834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  wt_actv_pvld_out_0_60 = _RAND_835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  wt_actv_pvld_out_0_61 = _RAND_836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  wt_actv_pvld_out_0_62 = _RAND_837[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  wt_actv_pvld_out_0_63 = _RAND_838[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  wt_actv_pvld_out_0_64 = _RAND_839[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  wt_actv_pvld_out_0_65 = _RAND_840[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  wt_actv_pvld_out_0_66 = _RAND_841[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  wt_actv_pvld_out_0_67 = _RAND_842[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  wt_actv_pvld_out_0_68 = _RAND_843[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  wt_actv_pvld_out_0_69 = _RAND_844[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  wt_actv_pvld_out_0_70 = _RAND_845[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  wt_actv_pvld_out_0_71 = _RAND_846[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  wt_actv_pvld_out_0_72 = _RAND_847[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  wt_actv_pvld_out_0_73 = _RAND_848[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  wt_actv_pvld_out_0_74 = _RAND_849[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  wt_actv_pvld_out_0_75 = _RAND_850[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  wt_actv_pvld_out_0_76 = _RAND_851[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  wt_actv_pvld_out_0_77 = _RAND_852[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  wt_actv_pvld_out_0_78 = _RAND_853[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  wt_actv_pvld_out_0_79 = _RAND_854[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  wt_actv_pvld_out_0_80 = _RAND_855[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  wt_actv_pvld_out_0_81 = _RAND_856[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  wt_actv_pvld_out_0_82 = _RAND_857[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  wt_actv_pvld_out_0_83 = _RAND_858[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  wt_actv_pvld_out_0_84 = _RAND_859[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  wt_actv_pvld_out_0_85 = _RAND_860[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  wt_actv_pvld_out_0_86 = _RAND_861[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  wt_actv_pvld_out_0_87 = _RAND_862[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  wt_actv_pvld_out_0_88 = _RAND_863[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  wt_actv_pvld_out_0_89 = _RAND_864[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  wt_actv_pvld_out_0_90 = _RAND_865[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  wt_actv_pvld_out_0_91 = _RAND_866[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  wt_actv_pvld_out_0_92 = _RAND_867[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  wt_actv_pvld_out_0_93 = _RAND_868[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  wt_actv_pvld_out_0_94 = _RAND_869[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  wt_actv_pvld_out_0_95 = _RAND_870[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  wt_actv_pvld_out_0_96 = _RAND_871[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  wt_actv_pvld_out_0_97 = _RAND_872[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  wt_actv_pvld_out_0_98 = _RAND_873[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  wt_actv_pvld_out_0_99 = _RAND_874[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  wt_actv_pvld_out_0_100 = _RAND_875[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  wt_actv_pvld_out_0_101 = _RAND_876[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  wt_actv_pvld_out_0_102 = _RAND_877[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  wt_actv_pvld_out_0_103 = _RAND_878[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  wt_actv_pvld_out_0_104 = _RAND_879[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  wt_actv_pvld_out_0_105 = _RAND_880[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  wt_actv_pvld_out_0_106 = _RAND_881[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  wt_actv_pvld_out_0_107 = _RAND_882[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  wt_actv_pvld_out_0_108 = _RAND_883[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  wt_actv_pvld_out_0_109 = _RAND_884[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  wt_actv_pvld_out_0_110 = _RAND_885[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  wt_actv_pvld_out_0_111 = _RAND_886[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  wt_actv_pvld_out_0_112 = _RAND_887[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  wt_actv_pvld_out_0_113 = _RAND_888[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  wt_actv_pvld_out_0_114 = _RAND_889[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  wt_actv_pvld_out_0_115 = _RAND_890[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  wt_actv_pvld_out_0_116 = _RAND_891[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  wt_actv_pvld_out_0_117 = _RAND_892[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  wt_actv_pvld_out_0_118 = _RAND_893[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  wt_actv_pvld_out_0_119 = _RAND_894[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  wt_actv_pvld_out_0_120 = _RAND_895[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  wt_actv_pvld_out_0_121 = _RAND_896[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  wt_actv_pvld_out_0_122 = _RAND_897[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  wt_actv_pvld_out_0_123 = _RAND_898[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  wt_actv_pvld_out_0_124 = _RAND_899[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  wt_actv_pvld_out_0_125 = _RAND_900[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  wt_actv_pvld_out_0_126 = _RAND_901[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  wt_actv_pvld_out_0_127 = _RAND_902[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  wt_actv_nz_out_0_0 = _RAND_903[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  wt_actv_nz_out_0_1 = _RAND_904[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  wt_actv_nz_out_0_2 = _RAND_905[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  wt_actv_nz_out_0_3 = _RAND_906[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  wt_actv_nz_out_0_4 = _RAND_907[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  wt_actv_nz_out_0_5 = _RAND_908[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  wt_actv_nz_out_0_6 = _RAND_909[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  wt_actv_nz_out_0_7 = _RAND_910[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  wt_actv_nz_out_0_8 = _RAND_911[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  wt_actv_nz_out_0_9 = _RAND_912[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  wt_actv_nz_out_0_10 = _RAND_913[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  wt_actv_nz_out_0_11 = _RAND_914[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  wt_actv_nz_out_0_12 = _RAND_915[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  wt_actv_nz_out_0_13 = _RAND_916[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  wt_actv_nz_out_0_14 = _RAND_917[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  wt_actv_nz_out_0_15 = _RAND_918[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  wt_actv_nz_out_0_16 = _RAND_919[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  wt_actv_nz_out_0_17 = _RAND_920[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  wt_actv_nz_out_0_18 = _RAND_921[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  wt_actv_nz_out_0_19 = _RAND_922[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  wt_actv_nz_out_0_20 = _RAND_923[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  wt_actv_nz_out_0_21 = _RAND_924[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  wt_actv_nz_out_0_22 = _RAND_925[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  wt_actv_nz_out_0_23 = _RAND_926[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  wt_actv_nz_out_0_24 = _RAND_927[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  wt_actv_nz_out_0_25 = _RAND_928[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  wt_actv_nz_out_0_26 = _RAND_929[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  wt_actv_nz_out_0_27 = _RAND_930[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  wt_actv_nz_out_0_28 = _RAND_931[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  wt_actv_nz_out_0_29 = _RAND_932[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  wt_actv_nz_out_0_30 = _RAND_933[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  wt_actv_nz_out_0_31 = _RAND_934[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  wt_actv_nz_out_0_32 = _RAND_935[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  wt_actv_nz_out_0_33 = _RAND_936[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  wt_actv_nz_out_0_34 = _RAND_937[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  wt_actv_nz_out_0_35 = _RAND_938[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  wt_actv_nz_out_0_36 = _RAND_939[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  wt_actv_nz_out_0_37 = _RAND_940[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  wt_actv_nz_out_0_38 = _RAND_941[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  wt_actv_nz_out_0_39 = _RAND_942[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  wt_actv_nz_out_0_40 = _RAND_943[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  wt_actv_nz_out_0_41 = _RAND_944[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  wt_actv_nz_out_0_42 = _RAND_945[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  wt_actv_nz_out_0_43 = _RAND_946[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  wt_actv_nz_out_0_44 = _RAND_947[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  wt_actv_nz_out_0_45 = _RAND_948[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  wt_actv_nz_out_0_46 = _RAND_949[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  wt_actv_nz_out_0_47 = _RAND_950[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  wt_actv_nz_out_0_48 = _RAND_951[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  wt_actv_nz_out_0_49 = _RAND_952[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  wt_actv_nz_out_0_50 = _RAND_953[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  wt_actv_nz_out_0_51 = _RAND_954[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  wt_actv_nz_out_0_52 = _RAND_955[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  wt_actv_nz_out_0_53 = _RAND_956[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  wt_actv_nz_out_0_54 = _RAND_957[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  wt_actv_nz_out_0_55 = _RAND_958[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  wt_actv_nz_out_0_56 = _RAND_959[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  wt_actv_nz_out_0_57 = _RAND_960[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  wt_actv_nz_out_0_58 = _RAND_961[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  wt_actv_nz_out_0_59 = _RAND_962[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  wt_actv_nz_out_0_60 = _RAND_963[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  wt_actv_nz_out_0_61 = _RAND_964[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  wt_actv_nz_out_0_62 = _RAND_965[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  wt_actv_nz_out_0_63 = _RAND_966[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  wt_actv_nz_out_0_64 = _RAND_967[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  wt_actv_nz_out_0_65 = _RAND_968[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  wt_actv_nz_out_0_66 = _RAND_969[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  wt_actv_nz_out_0_67 = _RAND_970[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  wt_actv_nz_out_0_68 = _RAND_971[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  wt_actv_nz_out_0_69 = _RAND_972[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  wt_actv_nz_out_0_70 = _RAND_973[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  wt_actv_nz_out_0_71 = _RAND_974[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  wt_actv_nz_out_0_72 = _RAND_975[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  wt_actv_nz_out_0_73 = _RAND_976[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  wt_actv_nz_out_0_74 = _RAND_977[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  wt_actv_nz_out_0_75 = _RAND_978[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  wt_actv_nz_out_0_76 = _RAND_979[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  wt_actv_nz_out_0_77 = _RAND_980[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  wt_actv_nz_out_0_78 = _RAND_981[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  wt_actv_nz_out_0_79 = _RAND_982[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  wt_actv_nz_out_0_80 = _RAND_983[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  wt_actv_nz_out_0_81 = _RAND_984[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  wt_actv_nz_out_0_82 = _RAND_985[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  wt_actv_nz_out_0_83 = _RAND_986[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  wt_actv_nz_out_0_84 = _RAND_987[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  wt_actv_nz_out_0_85 = _RAND_988[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  wt_actv_nz_out_0_86 = _RAND_989[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  wt_actv_nz_out_0_87 = _RAND_990[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  wt_actv_nz_out_0_88 = _RAND_991[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  wt_actv_nz_out_0_89 = _RAND_992[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  wt_actv_nz_out_0_90 = _RAND_993[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  wt_actv_nz_out_0_91 = _RAND_994[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  wt_actv_nz_out_0_92 = _RAND_995[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  wt_actv_nz_out_0_93 = _RAND_996[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  wt_actv_nz_out_0_94 = _RAND_997[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  wt_actv_nz_out_0_95 = _RAND_998[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  wt_actv_nz_out_0_96 = _RAND_999[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  wt_actv_nz_out_0_97 = _RAND_1000[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  wt_actv_nz_out_0_98 = _RAND_1001[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  wt_actv_nz_out_0_99 = _RAND_1002[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  wt_actv_nz_out_0_100 = _RAND_1003[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  wt_actv_nz_out_0_101 = _RAND_1004[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  wt_actv_nz_out_0_102 = _RAND_1005[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  wt_actv_nz_out_0_103 = _RAND_1006[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  wt_actv_nz_out_0_104 = _RAND_1007[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  wt_actv_nz_out_0_105 = _RAND_1008[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  wt_actv_nz_out_0_106 = _RAND_1009[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  wt_actv_nz_out_0_107 = _RAND_1010[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  wt_actv_nz_out_0_108 = _RAND_1011[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  wt_actv_nz_out_0_109 = _RAND_1012[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  wt_actv_nz_out_0_110 = _RAND_1013[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  wt_actv_nz_out_0_111 = _RAND_1014[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  wt_actv_nz_out_0_112 = _RAND_1015[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  wt_actv_nz_out_0_113 = _RAND_1016[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  wt_actv_nz_out_0_114 = _RAND_1017[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  wt_actv_nz_out_0_115 = _RAND_1018[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  wt_actv_nz_out_0_116 = _RAND_1019[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  wt_actv_nz_out_0_117 = _RAND_1020[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  wt_actv_nz_out_0_118 = _RAND_1021[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  wt_actv_nz_out_0_119 = _RAND_1022[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  wt_actv_nz_out_0_120 = _RAND_1023[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  wt_actv_nz_out_0_121 = _RAND_1024[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  wt_actv_nz_out_0_122 = _RAND_1025[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  wt_actv_nz_out_0_123 = _RAND_1026[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  wt_actv_nz_out_0_124 = _RAND_1027[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  wt_actv_nz_out_0_125 = _RAND_1028[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  wt_actv_nz_out_0_126 = _RAND_1029[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  wt_actv_nz_out_0_127 = _RAND_1030[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  wt_actv_data_out_0_0 = _RAND_1031[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  wt_actv_data_out_0_1 = _RAND_1032[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  wt_actv_data_out_0_2 = _RAND_1033[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  wt_actv_data_out_0_3 = _RAND_1034[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  wt_actv_data_out_0_4 = _RAND_1035[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  wt_actv_data_out_0_5 = _RAND_1036[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  wt_actv_data_out_0_6 = _RAND_1037[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  wt_actv_data_out_0_7 = _RAND_1038[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  wt_actv_data_out_0_8 = _RAND_1039[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  wt_actv_data_out_0_9 = _RAND_1040[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  wt_actv_data_out_0_10 = _RAND_1041[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  wt_actv_data_out_0_11 = _RAND_1042[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  wt_actv_data_out_0_12 = _RAND_1043[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  wt_actv_data_out_0_13 = _RAND_1044[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  wt_actv_data_out_0_14 = _RAND_1045[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  wt_actv_data_out_0_15 = _RAND_1046[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  wt_actv_data_out_0_16 = _RAND_1047[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  wt_actv_data_out_0_17 = _RAND_1048[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  wt_actv_data_out_0_18 = _RAND_1049[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  wt_actv_data_out_0_19 = _RAND_1050[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  wt_actv_data_out_0_20 = _RAND_1051[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  wt_actv_data_out_0_21 = _RAND_1052[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  wt_actv_data_out_0_22 = _RAND_1053[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  wt_actv_data_out_0_23 = _RAND_1054[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  wt_actv_data_out_0_24 = _RAND_1055[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  wt_actv_data_out_0_25 = _RAND_1056[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  wt_actv_data_out_0_26 = _RAND_1057[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  wt_actv_data_out_0_27 = _RAND_1058[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  wt_actv_data_out_0_28 = _RAND_1059[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  wt_actv_data_out_0_29 = _RAND_1060[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  wt_actv_data_out_0_30 = _RAND_1061[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  wt_actv_data_out_0_31 = _RAND_1062[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  wt_actv_data_out_0_32 = _RAND_1063[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  wt_actv_data_out_0_33 = _RAND_1064[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  wt_actv_data_out_0_34 = _RAND_1065[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  wt_actv_data_out_0_35 = _RAND_1066[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  wt_actv_data_out_0_36 = _RAND_1067[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  wt_actv_data_out_0_37 = _RAND_1068[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  wt_actv_data_out_0_38 = _RAND_1069[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  wt_actv_data_out_0_39 = _RAND_1070[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  wt_actv_data_out_0_40 = _RAND_1071[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  wt_actv_data_out_0_41 = _RAND_1072[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  wt_actv_data_out_0_42 = _RAND_1073[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  wt_actv_data_out_0_43 = _RAND_1074[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  wt_actv_data_out_0_44 = _RAND_1075[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  wt_actv_data_out_0_45 = _RAND_1076[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  wt_actv_data_out_0_46 = _RAND_1077[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  wt_actv_data_out_0_47 = _RAND_1078[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  wt_actv_data_out_0_48 = _RAND_1079[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  wt_actv_data_out_0_49 = _RAND_1080[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  wt_actv_data_out_0_50 = _RAND_1081[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  wt_actv_data_out_0_51 = _RAND_1082[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  wt_actv_data_out_0_52 = _RAND_1083[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  wt_actv_data_out_0_53 = _RAND_1084[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  wt_actv_data_out_0_54 = _RAND_1085[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  wt_actv_data_out_0_55 = _RAND_1086[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  wt_actv_data_out_0_56 = _RAND_1087[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  wt_actv_data_out_0_57 = _RAND_1088[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  wt_actv_data_out_0_58 = _RAND_1089[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  wt_actv_data_out_0_59 = _RAND_1090[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  wt_actv_data_out_0_60 = _RAND_1091[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  wt_actv_data_out_0_61 = _RAND_1092[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  wt_actv_data_out_0_62 = _RAND_1093[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  wt_actv_data_out_0_63 = _RAND_1094[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{`RANDOM}};
  wt_actv_data_out_0_64 = _RAND_1095[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{`RANDOM}};
  wt_actv_data_out_0_65 = _RAND_1096[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{`RANDOM}};
  wt_actv_data_out_0_66 = _RAND_1097[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{`RANDOM}};
  wt_actv_data_out_0_67 = _RAND_1098[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{`RANDOM}};
  wt_actv_data_out_0_68 = _RAND_1099[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{`RANDOM}};
  wt_actv_data_out_0_69 = _RAND_1100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{`RANDOM}};
  wt_actv_data_out_0_70 = _RAND_1101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{`RANDOM}};
  wt_actv_data_out_0_71 = _RAND_1102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{`RANDOM}};
  wt_actv_data_out_0_72 = _RAND_1103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{`RANDOM}};
  wt_actv_data_out_0_73 = _RAND_1104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{`RANDOM}};
  wt_actv_data_out_0_74 = _RAND_1105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{`RANDOM}};
  wt_actv_data_out_0_75 = _RAND_1106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{`RANDOM}};
  wt_actv_data_out_0_76 = _RAND_1107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{`RANDOM}};
  wt_actv_data_out_0_77 = _RAND_1108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{`RANDOM}};
  wt_actv_data_out_0_78 = _RAND_1109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{`RANDOM}};
  wt_actv_data_out_0_79 = _RAND_1110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{`RANDOM}};
  wt_actv_data_out_0_80 = _RAND_1111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{`RANDOM}};
  wt_actv_data_out_0_81 = _RAND_1112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{`RANDOM}};
  wt_actv_data_out_0_82 = _RAND_1113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{`RANDOM}};
  wt_actv_data_out_0_83 = _RAND_1114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{`RANDOM}};
  wt_actv_data_out_0_84 = _RAND_1115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{`RANDOM}};
  wt_actv_data_out_0_85 = _RAND_1116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{`RANDOM}};
  wt_actv_data_out_0_86 = _RAND_1117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{`RANDOM}};
  wt_actv_data_out_0_87 = _RAND_1118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{`RANDOM}};
  wt_actv_data_out_0_88 = _RAND_1119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{`RANDOM}};
  wt_actv_data_out_0_89 = _RAND_1120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{`RANDOM}};
  wt_actv_data_out_0_90 = _RAND_1121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{`RANDOM}};
  wt_actv_data_out_0_91 = _RAND_1122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{`RANDOM}};
  wt_actv_data_out_0_92 = _RAND_1123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{`RANDOM}};
  wt_actv_data_out_0_93 = _RAND_1124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{`RANDOM}};
  wt_actv_data_out_0_94 = _RAND_1125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{`RANDOM}};
  wt_actv_data_out_0_95 = _RAND_1126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{`RANDOM}};
  wt_actv_data_out_0_96 = _RAND_1127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{`RANDOM}};
  wt_actv_data_out_0_97 = _RAND_1128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{`RANDOM}};
  wt_actv_data_out_0_98 = _RAND_1129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{`RANDOM}};
  wt_actv_data_out_0_99 = _RAND_1130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{`RANDOM}};
  wt_actv_data_out_0_100 = _RAND_1131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{`RANDOM}};
  wt_actv_data_out_0_101 = _RAND_1132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{`RANDOM}};
  wt_actv_data_out_0_102 = _RAND_1133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{`RANDOM}};
  wt_actv_data_out_0_103 = _RAND_1134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{`RANDOM}};
  wt_actv_data_out_0_104 = _RAND_1135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{`RANDOM}};
  wt_actv_data_out_0_105 = _RAND_1136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{`RANDOM}};
  wt_actv_data_out_0_106 = _RAND_1137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{`RANDOM}};
  wt_actv_data_out_0_107 = _RAND_1138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{`RANDOM}};
  wt_actv_data_out_0_108 = _RAND_1139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{`RANDOM}};
  wt_actv_data_out_0_109 = _RAND_1140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{`RANDOM}};
  wt_actv_data_out_0_110 = _RAND_1141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{`RANDOM}};
  wt_actv_data_out_0_111 = _RAND_1142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{`RANDOM}};
  wt_actv_data_out_0_112 = _RAND_1143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{`RANDOM}};
  wt_actv_data_out_0_113 = _RAND_1144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{`RANDOM}};
  wt_actv_data_out_0_114 = _RAND_1145[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{`RANDOM}};
  wt_actv_data_out_0_115 = _RAND_1146[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{`RANDOM}};
  wt_actv_data_out_0_116 = _RAND_1147[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{`RANDOM}};
  wt_actv_data_out_0_117 = _RAND_1148[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{`RANDOM}};
  wt_actv_data_out_0_118 = _RAND_1149[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{`RANDOM}};
  wt_actv_data_out_0_119 = _RAND_1150[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{`RANDOM}};
  wt_actv_data_out_0_120 = _RAND_1151[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{`RANDOM}};
  wt_actv_data_out_0_121 = _RAND_1152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{`RANDOM}};
  wt_actv_data_out_0_122 = _RAND_1153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{`RANDOM}};
  wt_actv_data_out_0_123 = _RAND_1154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{`RANDOM}};
  wt_actv_data_out_0_124 = _RAND_1155[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{`RANDOM}};
  wt_actv_data_out_0_125 = _RAND_1156[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{`RANDOM}};
  wt_actv_data_out_0_126 = _RAND_1157[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{`RANDOM}};
  wt_actv_data_out_0_127 = _RAND_1158[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{`RANDOM}};
  dat_actv_data_reg_0_0 = _RAND_1159[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{`RANDOM}};
  dat_actv_data_reg_0_1 = _RAND_1160[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{`RANDOM}};
  dat_actv_data_reg_0_2 = _RAND_1161[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{`RANDOM}};
  dat_actv_data_reg_0_3 = _RAND_1162[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{`RANDOM}};
  dat_actv_data_reg_0_4 = _RAND_1163[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{`RANDOM}};
  dat_actv_data_reg_0_5 = _RAND_1164[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{`RANDOM}};
  dat_actv_data_reg_0_6 = _RAND_1165[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{`RANDOM}};
  dat_actv_data_reg_0_7 = _RAND_1166[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{`RANDOM}};
  dat_actv_data_reg_0_8 = _RAND_1167[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{`RANDOM}};
  dat_actv_data_reg_0_9 = _RAND_1168[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{`RANDOM}};
  dat_actv_data_reg_0_10 = _RAND_1169[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{`RANDOM}};
  dat_actv_data_reg_0_11 = _RAND_1170[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{`RANDOM}};
  dat_actv_data_reg_0_12 = _RAND_1171[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{`RANDOM}};
  dat_actv_data_reg_0_13 = _RAND_1172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{`RANDOM}};
  dat_actv_data_reg_0_14 = _RAND_1173[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{`RANDOM}};
  dat_actv_data_reg_0_15 = _RAND_1174[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{`RANDOM}};
  dat_actv_data_reg_0_16 = _RAND_1175[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{`RANDOM}};
  dat_actv_data_reg_0_17 = _RAND_1176[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{`RANDOM}};
  dat_actv_data_reg_0_18 = _RAND_1177[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{`RANDOM}};
  dat_actv_data_reg_0_19 = _RAND_1178[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{`RANDOM}};
  dat_actv_data_reg_0_20 = _RAND_1179[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{`RANDOM}};
  dat_actv_data_reg_0_21 = _RAND_1180[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{`RANDOM}};
  dat_actv_data_reg_0_22 = _RAND_1181[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{`RANDOM}};
  dat_actv_data_reg_0_23 = _RAND_1182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{`RANDOM}};
  dat_actv_data_reg_0_24 = _RAND_1183[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{`RANDOM}};
  dat_actv_data_reg_0_25 = _RAND_1184[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{`RANDOM}};
  dat_actv_data_reg_0_26 = _RAND_1185[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{`RANDOM}};
  dat_actv_data_reg_0_27 = _RAND_1186[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{`RANDOM}};
  dat_actv_data_reg_0_28 = _RAND_1187[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{`RANDOM}};
  dat_actv_data_reg_0_29 = _RAND_1188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{`RANDOM}};
  dat_actv_data_reg_0_30 = _RAND_1189[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{`RANDOM}};
  dat_actv_data_reg_0_31 = _RAND_1190[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{`RANDOM}};
  dat_actv_data_reg_0_32 = _RAND_1191[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{`RANDOM}};
  dat_actv_data_reg_0_33 = _RAND_1192[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{`RANDOM}};
  dat_actv_data_reg_0_34 = _RAND_1193[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{`RANDOM}};
  dat_actv_data_reg_0_35 = _RAND_1194[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{`RANDOM}};
  dat_actv_data_reg_0_36 = _RAND_1195[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{`RANDOM}};
  dat_actv_data_reg_0_37 = _RAND_1196[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{`RANDOM}};
  dat_actv_data_reg_0_38 = _RAND_1197[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{`RANDOM}};
  dat_actv_data_reg_0_39 = _RAND_1198[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{`RANDOM}};
  dat_actv_data_reg_0_40 = _RAND_1199[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{`RANDOM}};
  dat_actv_data_reg_0_41 = _RAND_1200[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{`RANDOM}};
  dat_actv_data_reg_0_42 = _RAND_1201[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{`RANDOM}};
  dat_actv_data_reg_0_43 = _RAND_1202[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{`RANDOM}};
  dat_actv_data_reg_0_44 = _RAND_1203[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{`RANDOM}};
  dat_actv_data_reg_0_45 = _RAND_1204[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{`RANDOM}};
  dat_actv_data_reg_0_46 = _RAND_1205[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{`RANDOM}};
  dat_actv_data_reg_0_47 = _RAND_1206[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{`RANDOM}};
  dat_actv_data_reg_0_48 = _RAND_1207[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{`RANDOM}};
  dat_actv_data_reg_0_49 = _RAND_1208[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{`RANDOM}};
  dat_actv_data_reg_0_50 = _RAND_1209[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{`RANDOM}};
  dat_actv_data_reg_0_51 = _RAND_1210[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{`RANDOM}};
  dat_actv_data_reg_0_52 = _RAND_1211[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{`RANDOM}};
  dat_actv_data_reg_0_53 = _RAND_1212[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{`RANDOM}};
  dat_actv_data_reg_0_54 = _RAND_1213[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{`RANDOM}};
  dat_actv_data_reg_0_55 = _RAND_1214[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{`RANDOM}};
  dat_actv_data_reg_0_56 = _RAND_1215[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{`RANDOM}};
  dat_actv_data_reg_0_57 = _RAND_1216[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{`RANDOM}};
  dat_actv_data_reg_0_58 = _RAND_1217[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{`RANDOM}};
  dat_actv_data_reg_0_59 = _RAND_1218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{`RANDOM}};
  dat_actv_data_reg_0_60 = _RAND_1219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{`RANDOM}};
  dat_actv_data_reg_0_61 = _RAND_1220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{`RANDOM}};
  dat_actv_data_reg_0_62 = _RAND_1221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{`RANDOM}};
  dat_actv_data_reg_0_63 = _RAND_1222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{`RANDOM}};
  dat_actv_data_reg_0_64 = _RAND_1223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{`RANDOM}};
  dat_actv_data_reg_0_65 = _RAND_1224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{`RANDOM}};
  dat_actv_data_reg_0_66 = _RAND_1225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{`RANDOM}};
  dat_actv_data_reg_0_67 = _RAND_1226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{`RANDOM}};
  dat_actv_data_reg_0_68 = _RAND_1227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{`RANDOM}};
  dat_actv_data_reg_0_69 = _RAND_1228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{`RANDOM}};
  dat_actv_data_reg_0_70 = _RAND_1229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{`RANDOM}};
  dat_actv_data_reg_0_71 = _RAND_1230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{`RANDOM}};
  dat_actv_data_reg_0_72 = _RAND_1231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{`RANDOM}};
  dat_actv_data_reg_0_73 = _RAND_1232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{`RANDOM}};
  dat_actv_data_reg_0_74 = _RAND_1233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{`RANDOM}};
  dat_actv_data_reg_0_75 = _RAND_1234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{`RANDOM}};
  dat_actv_data_reg_0_76 = _RAND_1235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{`RANDOM}};
  dat_actv_data_reg_0_77 = _RAND_1236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{`RANDOM}};
  dat_actv_data_reg_0_78 = _RAND_1237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{`RANDOM}};
  dat_actv_data_reg_0_79 = _RAND_1238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{`RANDOM}};
  dat_actv_data_reg_0_80 = _RAND_1239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{`RANDOM}};
  dat_actv_data_reg_0_81 = _RAND_1240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{`RANDOM}};
  dat_actv_data_reg_0_82 = _RAND_1241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{`RANDOM}};
  dat_actv_data_reg_0_83 = _RAND_1242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{`RANDOM}};
  dat_actv_data_reg_0_84 = _RAND_1243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{`RANDOM}};
  dat_actv_data_reg_0_85 = _RAND_1244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{`RANDOM}};
  dat_actv_data_reg_0_86 = _RAND_1245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{`RANDOM}};
  dat_actv_data_reg_0_87 = _RAND_1246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{`RANDOM}};
  dat_actv_data_reg_0_88 = _RAND_1247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{`RANDOM}};
  dat_actv_data_reg_0_89 = _RAND_1248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{`RANDOM}};
  dat_actv_data_reg_0_90 = _RAND_1249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{`RANDOM}};
  dat_actv_data_reg_0_91 = _RAND_1250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{`RANDOM}};
  dat_actv_data_reg_0_92 = _RAND_1251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1252 = {1{`RANDOM}};
  dat_actv_data_reg_0_93 = _RAND_1252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1253 = {1{`RANDOM}};
  dat_actv_data_reg_0_94 = _RAND_1253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1254 = {1{`RANDOM}};
  dat_actv_data_reg_0_95 = _RAND_1254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1255 = {1{`RANDOM}};
  dat_actv_data_reg_0_96 = _RAND_1255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1256 = {1{`RANDOM}};
  dat_actv_data_reg_0_97 = _RAND_1256[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1257 = {1{`RANDOM}};
  dat_actv_data_reg_0_98 = _RAND_1257[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1258 = {1{`RANDOM}};
  dat_actv_data_reg_0_99 = _RAND_1258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1259 = {1{`RANDOM}};
  dat_actv_data_reg_0_100 = _RAND_1259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1260 = {1{`RANDOM}};
  dat_actv_data_reg_0_101 = _RAND_1260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1261 = {1{`RANDOM}};
  dat_actv_data_reg_0_102 = _RAND_1261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1262 = {1{`RANDOM}};
  dat_actv_data_reg_0_103 = _RAND_1262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1263 = {1{`RANDOM}};
  dat_actv_data_reg_0_104 = _RAND_1263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1264 = {1{`RANDOM}};
  dat_actv_data_reg_0_105 = _RAND_1264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1265 = {1{`RANDOM}};
  dat_actv_data_reg_0_106 = _RAND_1265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1266 = {1{`RANDOM}};
  dat_actv_data_reg_0_107 = _RAND_1266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1267 = {1{`RANDOM}};
  dat_actv_data_reg_0_108 = _RAND_1267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1268 = {1{`RANDOM}};
  dat_actv_data_reg_0_109 = _RAND_1268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1269 = {1{`RANDOM}};
  dat_actv_data_reg_0_110 = _RAND_1269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1270 = {1{`RANDOM}};
  dat_actv_data_reg_0_111 = _RAND_1270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1271 = {1{`RANDOM}};
  dat_actv_data_reg_0_112 = _RAND_1271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1272 = {1{`RANDOM}};
  dat_actv_data_reg_0_113 = _RAND_1272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1273 = {1{`RANDOM}};
  dat_actv_data_reg_0_114 = _RAND_1273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1274 = {1{`RANDOM}};
  dat_actv_data_reg_0_115 = _RAND_1274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1275 = {1{`RANDOM}};
  dat_actv_data_reg_0_116 = _RAND_1275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1276 = {1{`RANDOM}};
  dat_actv_data_reg_0_117 = _RAND_1276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1277 = {1{`RANDOM}};
  dat_actv_data_reg_0_118 = _RAND_1277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1278 = {1{`RANDOM}};
  dat_actv_data_reg_0_119 = _RAND_1278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1279 = {1{`RANDOM}};
  dat_actv_data_reg_0_120 = _RAND_1279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1280 = {1{`RANDOM}};
  dat_actv_data_reg_0_121 = _RAND_1280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1281 = {1{`RANDOM}};
  dat_actv_data_reg_0_122 = _RAND_1281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1282 = {1{`RANDOM}};
  dat_actv_data_reg_0_123 = _RAND_1282[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1283 = {1{`RANDOM}};
  dat_actv_data_reg_0_124 = _RAND_1283[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1284 = {1{`RANDOM}};
  dat_actv_data_reg_0_125 = _RAND_1284[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1285 = {1{`RANDOM}};
  dat_actv_data_reg_0_126 = _RAND_1285[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1286 = {1{`RANDOM}};
  dat_actv_data_reg_0_127 = _RAND_1286[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1287 = {1{`RANDOM}};
  dat_actv_nz_reg_0_0 = _RAND_1287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1288 = {1{`RANDOM}};
  dat_actv_nz_reg_0_1 = _RAND_1288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1289 = {1{`RANDOM}};
  dat_actv_nz_reg_0_2 = _RAND_1289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1290 = {1{`RANDOM}};
  dat_actv_nz_reg_0_3 = _RAND_1290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1291 = {1{`RANDOM}};
  dat_actv_nz_reg_0_4 = _RAND_1291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1292 = {1{`RANDOM}};
  dat_actv_nz_reg_0_5 = _RAND_1292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1293 = {1{`RANDOM}};
  dat_actv_nz_reg_0_6 = _RAND_1293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1294 = {1{`RANDOM}};
  dat_actv_nz_reg_0_7 = _RAND_1294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1295 = {1{`RANDOM}};
  dat_actv_nz_reg_0_8 = _RAND_1295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1296 = {1{`RANDOM}};
  dat_actv_nz_reg_0_9 = _RAND_1296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1297 = {1{`RANDOM}};
  dat_actv_nz_reg_0_10 = _RAND_1297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1298 = {1{`RANDOM}};
  dat_actv_nz_reg_0_11 = _RAND_1298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1299 = {1{`RANDOM}};
  dat_actv_nz_reg_0_12 = _RAND_1299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1300 = {1{`RANDOM}};
  dat_actv_nz_reg_0_13 = _RAND_1300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1301 = {1{`RANDOM}};
  dat_actv_nz_reg_0_14 = _RAND_1301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1302 = {1{`RANDOM}};
  dat_actv_nz_reg_0_15 = _RAND_1302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1303 = {1{`RANDOM}};
  dat_actv_nz_reg_0_16 = _RAND_1303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1304 = {1{`RANDOM}};
  dat_actv_nz_reg_0_17 = _RAND_1304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1305 = {1{`RANDOM}};
  dat_actv_nz_reg_0_18 = _RAND_1305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1306 = {1{`RANDOM}};
  dat_actv_nz_reg_0_19 = _RAND_1306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1307 = {1{`RANDOM}};
  dat_actv_nz_reg_0_20 = _RAND_1307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1308 = {1{`RANDOM}};
  dat_actv_nz_reg_0_21 = _RAND_1308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1309 = {1{`RANDOM}};
  dat_actv_nz_reg_0_22 = _RAND_1309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1310 = {1{`RANDOM}};
  dat_actv_nz_reg_0_23 = _RAND_1310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1311 = {1{`RANDOM}};
  dat_actv_nz_reg_0_24 = _RAND_1311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1312 = {1{`RANDOM}};
  dat_actv_nz_reg_0_25 = _RAND_1312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1313 = {1{`RANDOM}};
  dat_actv_nz_reg_0_26 = _RAND_1313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1314 = {1{`RANDOM}};
  dat_actv_nz_reg_0_27 = _RAND_1314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1315 = {1{`RANDOM}};
  dat_actv_nz_reg_0_28 = _RAND_1315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1316 = {1{`RANDOM}};
  dat_actv_nz_reg_0_29 = _RAND_1316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1317 = {1{`RANDOM}};
  dat_actv_nz_reg_0_30 = _RAND_1317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1318 = {1{`RANDOM}};
  dat_actv_nz_reg_0_31 = _RAND_1318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1319 = {1{`RANDOM}};
  dat_actv_nz_reg_0_32 = _RAND_1319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1320 = {1{`RANDOM}};
  dat_actv_nz_reg_0_33 = _RAND_1320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1321 = {1{`RANDOM}};
  dat_actv_nz_reg_0_34 = _RAND_1321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1322 = {1{`RANDOM}};
  dat_actv_nz_reg_0_35 = _RAND_1322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1323 = {1{`RANDOM}};
  dat_actv_nz_reg_0_36 = _RAND_1323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1324 = {1{`RANDOM}};
  dat_actv_nz_reg_0_37 = _RAND_1324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1325 = {1{`RANDOM}};
  dat_actv_nz_reg_0_38 = _RAND_1325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1326 = {1{`RANDOM}};
  dat_actv_nz_reg_0_39 = _RAND_1326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1327 = {1{`RANDOM}};
  dat_actv_nz_reg_0_40 = _RAND_1327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1328 = {1{`RANDOM}};
  dat_actv_nz_reg_0_41 = _RAND_1328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1329 = {1{`RANDOM}};
  dat_actv_nz_reg_0_42 = _RAND_1329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1330 = {1{`RANDOM}};
  dat_actv_nz_reg_0_43 = _RAND_1330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1331 = {1{`RANDOM}};
  dat_actv_nz_reg_0_44 = _RAND_1331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1332 = {1{`RANDOM}};
  dat_actv_nz_reg_0_45 = _RAND_1332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1333 = {1{`RANDOM}};
  dat_actv_nz_reg_0_46 = _RAND_1333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1334 = {1{`RANDOM}};
  dat_actv_nz_reg_0_47 = _RAND_1334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1335 = {1{`RANDOM}};
  dat_actv_nz_reg_0_48 = _RAND_1335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1336 = {1{`RANDOM}};
  dat_actv_nz_reg_0_49 = _RAND_1336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1337 = {1{`RANDOM}};
  dat_actv_nz_reg_0_50 = _RAND_1337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1338 = {1{`RANDOM}};
  dat_actv_nz_reg_0_51 = _RAND_1338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1339 = {1{`RANDOM}};
  dat_actv_nz_reg_0_52 = _RAND_1339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1340 = {1{`RANDOM}};
  dat_actv_nz_reg_0_53 = _RAND_1340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1341 = {1{`RANDOM}};
  dat_actv_nz_reg_0_54 = _RAND_1341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1342 = {1{`RANDOM}};
  dat_actv_nz_reg_0_55 = _RAND_1342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1343 = {1{`RANDOM}};
  dat_actv_nz_reg_0_56 = _RAND_1343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1344 = {1{`RANDOM}};
  dat_actv_nz_reg_0_57 = _RAND_1344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1345 = {1{`RANDOM}};
  dat_actv_nz_reg_0_58 = _RAND_1345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1346 = {1{`RANDOM}};
  dat_actv_nz_reg_0_59 = _RAND_1346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1347 = {1{`RANDOM}};
  dat_actv_nz_reg_0_60 = _RAND_1347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1348 = {1{`RANDOM}};
  dat_actv_nz_reg_0_61 = _RAND_1348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1349 = {1{`RANDOM}};
  dat_actv_nz_reg_0_62 = _RAND_1349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1350 = {1{`RANDOM}};
  dat_actv_nz_reg_0_63 = _RAND_1350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1351 = {1{`RANDOM}};
  dat_actv_nz_reg_0_64 = _RAND_1351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1352 = {1{`RANDOM}};
  dat_actv_nz_reg_0_65 = _RAND_1352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1353 = {1{`RANDOM}};
  dat_actv_nz_reg_0_66 = _RAND_1353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1354 = {1{`RANDOM}};
  dat_actv_nz_reg_0_67 = _RAND_1354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1355 = {1{`RANDOM}};
  dat_actv_nz_reg_0_68 = _RAND_1355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1356 = {1{`RANDOM}};
  dat_actv_nz_reg_0_69 = _RAND_1356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1357 = {1{`RANDOM}};
  dat_actv_nz_reg_0_70 = _RAND_1357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1358 = {1{`RANDOM}};
  dat_actv_nz_reg_0_71 = _RAND_1358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1359 = {1{`RANDOM}};
  dat_actv_nz_reg_0_72 = _RAND_1359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1360 = {1{`RANDOM}};
  dat_actv_nz_reg_0_73 = _RAND_1360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1361 = {1{`RANDOM}};
  dat_actv_nz_reg_0_74 = _RAND_1361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1362 = {1{`RANDOM}};
  dat_actv_nz_reg_0_75 = _RAND_1362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1363 = {1{`RANDOM}};
  dat_actv_nz_reg_0_76 = _RAND_1363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1364 = {1{`RANDOM}};
  dat_actv_nz_reg_0_77 = _RAND_1364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1365 = {1{`RANDOM}};
  dat_actv_nz_reg_0_78 = _RAND_1365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1366 = {1{`RANDOM}};
  dat_actv_nz_reg_0_79 = _RAND_1366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1367 = {1{`RANDOM}};
  dat_actv_nz_reg_0_80 = _RAND_1367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1368 = {1{`RANDOM}};
  dat_actv_nz_reg_0_81 = _RAND_1368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1369 = {1{`RANDOM}};
  dat_actv_nz_reg_0_82 = _RAND_1369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1370 = {1{`RANDOM}};
  dat_actv_nz_reg_0_83 = _RAND_1370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1371 = {1{`RANDOM}};
  dat_actv_nz_reg_0_84 = _RAND_1371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1372 = {1{`RANDOM}};
  dat_actv_nz_reg_0_85 = _RAND_1372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1373 = {1{`RANDOM}};
  dat_actv_nz_reg_0_86 = _RAND_1373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1374 = {1{`RANDOM}};
  dat_actv_nz_reg_0_87 = _RAND_1374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1375 = {1{`RANDOM}};
  dat_actv_nz_reg_0_88 = _RAND_1375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1376 = {1{`RANDOM}};
  dat_actv_nz_reg_0_89 = _RAND_1376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1377 = {1{`RANDOM}};
  dat_actv_nz_reg_0_90 = _RAND_1377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1378 = {1{`RANDOM}};
  dat_actv_nz_reg_0_91 = _RAND_1378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1379 = {1{`RANDOM}};
  dat_actv_nz_reg_0_92 = _RAND_1379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1380 = {1{`RANDOM}};
  dat_actv_nz_reg_0_93 = _RAND_1380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1381 = {1{`RANDOM}};
  dat_actv_nz_reg_0_94 = _RAND_1381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1382 = {1{`RANDOM}};
  dat_actv_nz_reg_0_95 = _RAND_1382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1383 = {1{`RANDOM}};
  dat_actv_nz_reg_0_96 = _RAND_1383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1384 = {1{`RANDOM}};
  dat_actv_nz_reg_0_97 = _RAND_1384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1385 = {1{`RANDOM}};
  dat_actv_nz_reg_0_98 = _RAND_1385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1386 = {1{`RANDOM}};
  dat_actv_nz_reg_0_99 = _RAND_1386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1387 = {1{`RANDOM}};
  dat_actv_nz_reg_0_100 = _RAND_1387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1388 = {1{`RANDOM}};
  dat_actv_nz_reg_0_101 = _RAND_1388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1389 = {1{`RANDOM}};
  dat_actv_nz_reg_0_102 = _RAND_1389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1390 = {1{`RANDOM}};
  dat_actv_nz_reg_0_103 = _RAND_1390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1391 = {1{`RANDOM}};
  dat_actv_nz_reg_0_104 = _RAND_1391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1392 = {1{`RANDOM}};
  dat_actv_nz_reg_0_105 = _RAND_1392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1393 = {1{`RANDOM}};
  dat_actv_nz_reg_0_106 = _RAND_1393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1394 = {1{`RANDOM}};
  dat_actv_nz_reg_0_107 = _RAND_1394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1395 = {1{`RANDOM}};
  dat_actv_nz_reg_0_108 = _RAND_1395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1396 = {1{`RANDOM}};
  dat_actv_nz_reg_0_109 = _RAND_1396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1397 = {1{`RANDOM}};
  dat_actv_nz_reg_0_110 = _RAND_1397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1398 = {1{`RANDOM}};
  dat_actv_nz_reg_0_111 = _RAND_1398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1399 = {1{`RANDOM}};
  dat_actv_nz_reg_0_112 = _RAND_1399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1400 = {1{`RANDOM}};
  dat_actv_nz_reg_0_113 = _RAND_1400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1401 = {1{`RANDOM}};
  dat_actv_nz_reg_0_114 = _RAND_1401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1402 = {1{`RANDOM}};
  dat_actv_nz_reg_0_115 = _RAND_1402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1403 = {1{`RANDOM}};
  dat_actv_nz_reg_0_116 = _RAND_1403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1404 = {1{`RANDOM}};
  dat_actv_nz_reg_0_117 = _RAND_1404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1405 = {1{`RANDOM}};
  dat_actv_nz_reg_0_118 = _RAND_1405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1406 = {1{`RANDOM}};
  dat_actv_nz_reg_0_119 = _RAND_1406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1407 = {1{`RANDOM}};
  dat_actv_nz_reg_0_120 = _RAND_1407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1408 = {1{`RANDOM}};
  dat_actv_nz_reg_0_121 = _RAND_1408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1409 = {1{`RANDOM}};
  dat_actv_nz_reg_0_122 = _RAND_1409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1410 = {1{`RANDOM}};
  dat_actv_nz_reg_0_123 = _RAND_1410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1411 = {1{`RANDOM}};
  dat_actv_nz_reg_0_124 = _RAND_1411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1412 = {1{`RANDOM}};
  dat_actv_nz_reg_0_125 = _RAND_1412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1413 = {1{`RANDOM}};
  dat_actv_nz_reg_0_126 = _RAND_1413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1414 = {1{`RANDOM}};
  dat_actv_nz_reg_0_127 = _RAND_1414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1415 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_0 = _RAND_1415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1416 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_1 = _RAND_1416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1417 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_2 = _RAND_1417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1418 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_3 = _RAND_1418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1419 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_4 = _RAND_1419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1420 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_5 = _RAND_1420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1421 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_6 = _RAND_1421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1422 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_7 = _RAND_1422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1423 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_8 = _RAND_1423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1424 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_9 = _RAND_1424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1425 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_10 = _RAND_1425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1426 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_11 = _RAND_1426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1427 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_12 = _RAND_1427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1428 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_13 = _RAND_1428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1429 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_14 = _RAND_1429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1430 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_15 = _RAND_1430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1431 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_16 = _RAND_1431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1432 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_17 = _RAND_1432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1433 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_18 = _RAND_1433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1434 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_19 = _RAND_1434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1435 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_20 = _RAND_1435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1436 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_21 = _RAND_1436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1437 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_22 = _RAND_1437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1438 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_23 = _RAND_1438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1439 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_24 = _RAND_1439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1440 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_25 = _RAND_1440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1441 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_26 = _RAND_1441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1442 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_27 = _RAND_1442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1443 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_28 = _RAND_1443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1444 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_29 = _RAND_1444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1445 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_30 = _RAND_1445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1446 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_31 = _RAND_1446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1447 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_32 = _RAND_1447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1448 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_33 = _RAND_1448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1449 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_34 = _RAND_1449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1450 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_35 = _RAND_1450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1451 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_36 = _RAND_1451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1452 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_37 = _RAND_1452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1453 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_38 = _RAND_1453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1454 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_39 = _RAND_1454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1455 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_40 = _RAND_1455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1456 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_41 = _RAND_1456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1457 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_42 = _RAND_1457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1458 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_43 = _RAND_1458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1459 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_44 = _RAND_1459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1460 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_45 = _RAND_1460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1461 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_46 = _RAND_1461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1462 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_47 = _RAND_1462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1463 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_48 = _RAND_1463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1464 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_49 = _RAND_1464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1465 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_50 = _RAND_1465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1466 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_51 = _RAND_1466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1467 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_52 = _RAND_1467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1468 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_53 = _RAND_1468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1469 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_54 = _RAND_1469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1470 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_55 = _RAND_1470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1471 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_56 = _RAND_1471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1472 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_57 = _RAND_1472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1473 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_58 = _RAND_1473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1474 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_59 = _RAND_1474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1475 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_60 = _RAND_1475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1476 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_61 = _RAND_1476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1477 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_62 = _RAND_1477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1478 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_63 = _RAND_1478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1479 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_64 = _RAND_1479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1480 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_65 = _RAND_1480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1481 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_66 = _RAND_1481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1482 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_67 = _RAND_1482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1483 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_68 = _RAND_1483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1484 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_69 = _RAND_1484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1485 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_70 = _RAND_1485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1486 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_71 = _RAND_1486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1487 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_72 = _RAND_1487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1488 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_73 = _RAND_1488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1489 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_74 = _RAND_1489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1490 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_75 = _RAND_1490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1491 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_76 = _RAND_1491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1492 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_77 = _RAND_1492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1493 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_78 = _RAND_1493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1494 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_79 = _RAND_1494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1495 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_80 = _RAND_1495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1496 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_81 = _RAND_1496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1497 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_82 = _RAND_1497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1498 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_83 = _RAND_1498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1499 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_84 = _RAND_1499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1500 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_85 = _RAND_1500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1501 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_86 = _RAND_1501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1502 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_87 = _RAND_1502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1503 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_88 = _RAND_1503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1504 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_89 = _RAND_1504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1505 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_90 = _RAND_1505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1506 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_91 = _RAND_1506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1507 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_92 = _RAND_1507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1508 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_93 = _RAND_1508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1509 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_94 = _RAND_1509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1510 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_95 = _RAND_1510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1511 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_96 = _RAND_1511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1512 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_97 = _RAND_1512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1513 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_98 = _RAND_1513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1514 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_99 = _RAND_1514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1515 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_100 = _RAND_1515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1516 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_101 = _RAND_1516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1517 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_102 = _RAND_1517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1518 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_103 = _RAND_1518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1519 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_104 = _RAND_1519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1520 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_105 = _RAND_1520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1521 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_106 = _RAND_1521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1522 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_107 = _RAND_1522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1523 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_108 = _RAND_1523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1524 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_109 = _RAND_1524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1525 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_110 = _RAND_1525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1526 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_111 = _RAND_1526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1527 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_112 = _RAND_1527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1528 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_113 = _RAND_1528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1529 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_114 = _RAND_1529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1530 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_115 = _RAND_1530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1531 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_116 = _RAND_1531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1532 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_117 = _RAND_1532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1533 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_118 = _RAND_1533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1534 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_119 = _RAND_1534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1535 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_120 = _RAND_1535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1536 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_121 = _RAND_1536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1537 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_122 = _RAND_1537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1538 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_123 = _RAND_1538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1539 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_124 = _RAND_1539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1540 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_125 = _RAND_1540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1541 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_126 = _RAND_1541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1542 = {1{`RANDOM}};
  dat_actv_pvld_reg_0_127 = _RAND_1542[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wt_pre_nz_0 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_0 <= io_in_wt_mask_0;
      end
    end
    if (reset) begin
      wt_pre_nz_1 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_1 <= io_in_wt_mask_1;
      end
    end
    if (reset) begin
      wt_pre_nz_2 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_2 <= io_in_wt_mask_2;
      end
    end
    if (reset) begin
      wt_pre_nz_3 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_3 <= io_in_wt_mask_3;
      end
    end
    if (reset) begin
      wt_pre_nz_4 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_4 <= io_in_wt_mask_4;
      end
    end
    if (reset) begin
      wt_pre_nz_5 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_5 <= io_in_wt_mask_5;
      end
    end
    if (reset) begin
      wt_pre_nz_6 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_6 <= io_in_wt_mask_6;
      end
    end
    if (reset) begin
      wt_pre_nz_7 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_7 <= io_in_wt_mask_7;
      end
    end
    if (reset) begin
      wt_pre_nz_8 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_8 <= io_in_wt_mask_8;
      end
    end
    if (reset) begin
      wt_pre_nz_9 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_9 <= io_in_wt_mask_9;
      end
    end
    if (reset) begin
      wt_pre_nz_10 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_10 <= io_in_wt_mask_10;
      end
    end
    if (reset) begin
      wt_pre_nz_11 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_11 <= io_in_wt_mask_11;
      end
    end
    if (reset) begin
      wt_pre_nz_12 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_12 <= io_in_wt_mask_12;
      end
    end
    if (reset) begin
      wt_pre_nz_13 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_13 <= io_in_wt_mask_13;
      end
    end
    if (reset) begin
      wt_pre_nz_14 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_14 <= io_in_wt_mask_14;
      end
    end
    if (reset) begin
      wt_pre_nz_15 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_15 <= io_in_wt_mask_15;
      end
    end
    if (reset) begin
      wt_pre_nz_16 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_16 <= io_in_wt_mask_16;
      end
    end
    if (reset) begin
      wt_pre_nz_17 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_17 <= io_in_wt_mask_17;
      end
    end
    if (reset) begin
      wt_pre_nz_18 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_18 <= io_in_wt_mask_18;
      end
    end
    if (reset) begin
      wt_pre_nz_19 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_19 <= io_in_wt_mask_19;
      end
    end
    if (reset) begin
      wt_pre_nz_20 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_20 <= io_in_wt_mask_20;
      end
    end
    if (reset) begin
      wt_pre_nz_21 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_21 <= io_in_wt_mask_21;
      end
    end
    if (reset) begin
      wt_pre_nz_22 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_22 <= io_in_wt_mask_22;
      end
    end
    if (reset) begin
      wt_pre_nz_23 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_23 <= io_in_wt_mask_23;
      end
    end
    if (reset) begin
      wt_pre_nz_24 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_24 <= io_in_wt_mask_24;
      end
    end
    if (reset) begin
      wt_pre_nz_25 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_25 <= io_in_wt_mask_25;
      end
    end
    if (reset) begin
      wt_pre_nz_26 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_26 <= io_in_wt_mask_26;
      end
    end
    if (reset) begin
      wt_pre_nz_27 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_27 <= io_in_wt_mask_27;
      end
    end
    if (reset) begin
      wt_pre_nz_28 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_28 <= io_in_wt_mask_28;
      end
    end
    if (reset) begin
      wt_pre_nz_29 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_29 <= io_in_wt_mask_29;
      end
    end
    if (reset) begin
      wt_pre_nz_30 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_30 <= io_in_wt_mask_30;
      end
    end
    if (reset) begin
      wt_pre_nz_31 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_31 <= io_in_wt_mask_31;
      end
    end
    if (reset) begin
      wt_pre_nz_32 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_32 <= io_in_wt_mask_32;
      end
    end
    if (reset) begin
      wt_pre_nz_33 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_33 <= io_in_wt_mask_33;
      end
    end
    if (reset) begin
      wt_pre_nz_34 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_34 <= io_in_wt_mask_34;
      end
    end
    if (reset) begin
      wt_pre_nz_35 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_35 <= io_in_wt_mask_35;
      end
    end
    if (reset) begin
      wt_pre_nz_36 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_36 <= io_in_wt_mask_36;
      end
    end
    if (reset) begin
      wt_pre_nz_37 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_37 <= io_in_wt_mask_37;
      end
    end
    if (reset) begin
      wt_pre_nz_38 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_38 <= io_in_wt_mask_38;
      end
    end
    if (reset) begin
      wt_pre_nz_39 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_39 <= io_in_wt_mask_39;
      end
    end
    if (reset) begin
      wt_pre_nz_40 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_40 <= io_in_wt_mask_40;
      end
    end
    if (reset) begin
      wt_pre_nz_41 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_41 <= io_in_wt_mask_41;
      end
    end
    if (reset) begin
      wt_pre_nz_42 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_42 <= io_in_wt_mask_42;
      end
    end
    if (reset) begin
      wt_pre_nz_43 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_43 <= io_in_wt_mask_43;
      end
    end
    if (reset) begin
      wt_pre_nz_44 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_44 <= io_in_wt_mask_44;
      end
    end
    if (reset) begin
      wt_pre_nz_45 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_45 <= io_in_wt_mask_45;
      end
    end
    if (reset) begin
      wt_pre_nz_46 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_46 <= io_in_wt_mask_46;
      end
    end
    if (reset) begin
      wt_pre_nz_47 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_47 <= io_in_wt_mask_47;
      end
    end
    if (reset) begin
      wt_pre_nz_48 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_48 <= io_in_wt_mask_48;
      end
    end
    if (reset) begin
      wt_pre_nz_49 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_49 <= io_in_wt_mask_49;
      end
    end
    if (reset) begin
      wt_pre_nz_50 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_50 <= io_in_wt_mask_50;
      end
    end
    if (reset) begin
      wt_pre_nz_51 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_51 <= io_in_wt_mask_51;
      end
    end
    if (reset) begin
      wt_pre_nz_52 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_52 <= io_in_wt_mask_52;
      end
    end
    if (reset) begin
      wt_pre_nz_53 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_53 <= io_in_wt_mask_53;
      end
    end
    if (reset) begin
      wt_pre_nz_54 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_54 <= io_in_wt_mask_54;
      end
    end
    if (reset) begin
      wt_pre_nz_55 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_55 <= io_in_wt_mask_55;
      end
    end
    if (reset) begin
      wt_pre_nz_56 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_56 <= io_in_wt_mask_56;
      end
    end
    if (reset) begin
      wt_pre_nz_57 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_57 <= io_in_wt_mask_57;
      end
    end
    if (reset) begin
      wt_pre_nz_58 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_58 <= io_in_wt_mask_58;
      end
    end
    if (reset) begin
      wt_pre_nz_59 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_59 <= io_in_wt_mask_59;
      end
    end
    if (reset) begin
      wt_pre_nz_60 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_60 <= io_in_wt_mask_60;
      end
    end
    if (reset) begin
      wt_pre_nz_61 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_61 <= io_in_wt_mask_61;
      end
    end
    if (reset) begin
      wt_pre_nz_62 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_62 <= io_in_wt_mask_62;
      end
    end
    if (reset) begin
      wt_pre_nz_63 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_63 <= io_in_wt_mask_63;
      end
    end
    if (reset) begin
      wt_pre_nz_64 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_64 <= io_in_wt_mask_64;
      end
    end
    if (reset) begin
      wt_pre_nz_65 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_65 <= io_in_wt_mask_65;
      end
    end
    if (reset) begin
      wt_pre_nz_66 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_66 <= io_in_wt_mask_66;
      end
    end
    if (reset) begin
      wt_pre_nz_67 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_67 <= io_in_wt_mask_67;
      end
    end
    if (reset) begin
      wt_pre_nz_68 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_68 <= io_in_wt_mask_68;
      end
    end
    if (reset) begin
      wt_pre_nz_69 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_69 <= io_in_wt_mask_69;
      end
    end
    if (reset) begin
      wt_pre_nz_70 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_70 <= io_in_wt_mask_70;
      end
    end
    if (reset) begin
      wt_pre_nz_71 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_71 <= io_in_wt_mask_71;
      end
    end
    if (reset) begin
      wt_pre_nz_72 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_72 <= io_in_wt_mask_72;
      end
    end
    if (reset) begin
      wt_pre_nz_73 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_73 <= io_in_wt_mask_73;
      end
    end
    if (reset) begin
      wt_pre_nz_74 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_74 <= io_in_wt_mask_74;
      end
    end
    if (reset) begin
      wt_pre_nz_75 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_75 <= io_in_wt_mask_75;
      end
    end
    if (reset) begin
      wt_pre_nz_76 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_76 <= io_in_wt_mask_76;
      end
    end
    if (reset) begin
      wt_pre_nz_77 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_77 <= io_in_wt_mask_77;
      end
    end
    if (reset) begin
      wt_pre_nz_78 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_78 <= io_in_wt_mask_78;
      end
    end
    if (reset) begin
      wt_pre_nz_79 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_79 <= io_in_wt_mask_79;
      end
    end
    if (reset) begin
      wt_pre_nz_80 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_80 <= io_in_wt_mask_80;
      end
    end
    if (reset) begin
      wt_pre_nz_81 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_81 <= io_in_wt_mask_81;
      end
    end
    if (reset) begin
      wt_pre_nz_82 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_82 <= io_in_wt_mask_82;
      end
    end
    if (reset) begin
      wt_pre_nz_83 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_83 <= io_in_wt_mask_83;
      end
    end
    if (reset) begin
      wt_pre_nz_84 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_84 <= io_in_wt_mask_84;
      end
    end
    if (reset) begin
      wt_pre_nz_85 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_85 <= io_in_wt_mask_85;
      end
    end
    if (reset) begin
      wt_pre_nz_86 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_86 <= io_in_wt_mask_86;
      end
    end
    if (reset) begin
      wt_pre_nz_87 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_87 <= io_in_wt_mask_87;
      end
    end
    if (reset) begin
      wt_pre_nz_88 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_88 <= io_in_wt_mask_88;
      end
    end
    if (reset) begin
      wt_pre_nz_89 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_89 <= io_in_wt_mask_89;
      end
    end
    if (reset) begin
      wt_pre_nz_90 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_90 <= io_in_wt_mask_90;
      end
    end
    if (reset) begin
      wt_pre_nz_91 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_91 <= io_in_wt_mask_91;
      end
    end
    if (reset) begin
      wt_pre_nz_92 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_92 <= io_in_wt_mask_92;
      end
    end
    if (reset) begin
      wt_pre_nz_93 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_93 <= io_in_wt_mask_93;
      end
    end
    if (reset) begin
      wt_pre_nz_94 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_94 <= io_in_wt_mask_94;
      end
    end
    if (reset) begin
      wt_pre_nz_95 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_95 <= io_in_wt_mask_95;
      end
    end
    if (reset) begin
      wt_pre_nz_96 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_96 <= io_in_wt_mask_96;
      end
    end
    if (reset) begin
      wt_pre_nz_97 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_97 <= io_in_wt_mask_97;
      end
    end
    if (reset) begin
      wt_pre_nz_98 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_98 <= io_in_wt_mask_98;
      end
    end
    if (reset) begin
      wt_pre_nz_99 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_99 <= io_in_wt_mask_99;
      end
    end
    if (reset) begin
      wt_pre_nz_100 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_100 <= io_in_wt_mask_100;
      end
    end
    if (reset) begin
      wt_pre_nz_101 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_101 <= io_in_wt_mask_101;
      end
    end
    if (reset) begin
      wt_pre_nz_102 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_102 <= io_in_wt_mask_102;
      end
    end
    if (reset) begin
      wt_pre_nz_103 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_103 <= io_in_wt_mask_103;
      end
    end
    if (reset) begin
      wt_pre_nz_104 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_104 <= io_in_wt_mask_104;
      end
    end
    if (reset) begin
      wt_pre_nz_105 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_105 <= io_in_wt_mask_105;
      end
    end
    if (reset) begin
      wt_pre_nz_106 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_106 <= io_in_wt_mask_106;
      end
    end
    if (reset) begin
      wt_pre_nz_107 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_107 <= io_in_wt_mask_107;
      end
    end
    if (reset) begin
      wt_pre_nz_108 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_108 <= io_in_wt_mask_108;
      end
    end
    if (reset) begin
      wt_pre_nz_109 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_109 <= io_in_wt_mask_109;
      end
    end
    if (reset) begin
      wt_pre_nz_110 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_110 <= io_in_wt_mask_110;
      end
    end
    if (reset) begin
      wt_pre_nz_111 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_111 <= io_in_wt_mask_111;
      end
    end
    if (reset) begin
      wt_pre_nz_112 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_112 <= io_in_wt_mask_112;
      end
    end
    if (reset) begin
      wt_pre_nz_113 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_113 <= io_in_wt_mask_113;
      end
    end
    if (reset) begin
      wt_pre_nz_114 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_114 <= io_in_wt_mask_114;
      end
    end
    if (reset) begin
      wt_pre_nz_115 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_115 <= io_in_wt_mask_115;
      end
    end
    if (reset) begin
      wt_pre_nz_116 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_116 <= io_in_wt_mask_116;
      end
    end
    if (reset) begin
      wt_pre_nz_117 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_117 <= io_in_wt_mask_117;
      end
    end
    if (reset) begin
      wt_pre_nz_118 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_118 <= io_in_wt_mask_118;
      end
    end
    if (reset) begin
      wt_pre_nz_119 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_119 <= io_in_wt_mask_119;
      end
    end
    if (reset) begin
      wt_pre_nz_120 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_120 <= io_in_wt_mask_120;
      end
    end
    if (reset) begin
      wt_pre_nz_121 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_121 <= io_in_wt_mask_121;
      end
    end
    if (reset) begin
      wt_pre_nz_122 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_122 <= io_in_wt_mask_122;
      end
    end
    if (reset) begin
      wt_pre_nz_123 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_123 <= io_in_wt_mask_123;
      end
    end
    if (reset) begin
      wt_pre_nz_124 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_124 <= io_in_wt_mask_124;
      end
    end
    if (reset) begin
      wt_pre_nz_125 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_125 <= io_in_wt_mask_125;
      end
    end
    if (reset) begin
      wt_pre_nz_126 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_126 <= io_in_wt_mask_126;
      end
    end
    if (reset) begin
      wt_pre_nz_127 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_nz_127 <= io_in_wt_mask_127;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_0) begin
        wt_pre_data_0 <= io_in_wt_data_0;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_1) begin
        wt_pre_data_1 <= io_in_wt_data_1;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_2) begin
        wt_pre_data_2 <= io_in_wt_data_2;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_3) begin
        wt_pre_data_3 <= io_in_wt_data_3;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_4) begin
        wt_pre_data_4 <= io_in_wt_data_4;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_5) begin
        wt_pre_data_5 <= io_in_wt_data_5;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_6) begin
        wt_pre_data_6 <= io_in_wt_data_6;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_7) begin
        wt_pre_data_7 <= io_in_wt_data_7;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_8) begin
        wt_pre_data_8 <= io_in_wt_data_8;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_9) begin
        wt_pre_data_9 <= io_in_wt_data_9;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_10) begin
        wt_pre_data_10 <= io_in_wt_data_10;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_11) begin
        wt_pre_data_11 <= io_in_wt_data_11;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_12) begin
        wt_pre_data_12 <= io_in_wt_data_12;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_13) begin
        wt_pre_data_13 <= io_in_wt_data_13;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_14) begin
        wt_pre_data_14 <= io_in_wt_data_14;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_15) begin
        wt_pre_data_15 <= io_in_wt_data_15;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_16) begin
        wt_pre_data_16 <= io_in_wt_data_16;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_17) begin
        wt_pre_data_17 <= io_in_wt_data_17;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_18) begin
        wt_pre_data_18 <= io_in_wt_data_18;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_19) begin
        wt_pre_data_19 <= io_in_wt_data_19;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_20) begin
        wt_pre_data_20 <= io_in_wt_data_20;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_21) begin
        wt_pre_data_21 <= io_in_wt_data_21;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_22) begin
        wt_pre_data_22 <= io_in_wt_data_22;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_23) begin
        wt_pre_data_23 <= io_in_wt_data_23;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_24) begin
        wt_pre_data_24 <= io_in_wt_data_24;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_25) begin
        wt_pre_data_25 <= io_in_wt_data_25;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_26) begin
        wt_pre_data_26 <= io_in_wt_data_26;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_27) begin
        wt_pre_data_27 <= io_in_wt_data_27;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_28) begin
        wt_pre_data_28 <= io_in_wt_data_28;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_29) begin
        wt_pre_data_29 <= io_in_wt_data_29;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_30) begin
        wt_pre_data_30 <= io_in_wt_data_30;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_31) begin
        wt_pre_data_31 <= io_in_wt_data_31;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_32) begin
        wt_pre_data_32 <= io_in_wt_data_32;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_33) begin
        wt_pre_data_33 <= io_in_wt_data_33;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_34) begin
        wt_pre_data_34 <= io_in_wt_data_34;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_35) begin
        wt_pre_data_35 <= io_in_wt_data_35;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_36) begin
        wt_pre_data_36 <= io_in_wt_data_36;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_37) begin
        wt_pre_data_37 <= io_in_wt_data_37;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_38) begin
        wt_pre_data_38 <= io_in_wt_data_38;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_39) begin
        wt_pre_data_39 <= io_in_wt_data_39;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_40) begin
        wt_pre_data_40 <= io_in_wt_data_40;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_41) begin
        wt_pre_data_41 <= io_in_wt_data_41;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_42) begin
        wt_pre_data_42 <= io_in_wt_data_42;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_43) begin
        wt_pre_data_43 <= io_in_wt_data_43;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_44) begin
        wt_pre_data_44 <= io_in_wt_data_44;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_45) begin
        wt_pre_data_45 <= io_in_wt_data_45;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_46) begin
        wt_pre_data_46 <= io_in_wt_data_46;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_47) begin
        wt_pre_data_47 <= io_in_wt_data_47;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_48) begin
        wt_pre_data_48 <= io_in_wt_data_48;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_49) begin
        wt_pre_data_49 <= io_in_wt_data_49;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_50) begin
        wt_pre_data_50 <= io_in_wt_data_50;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_51) begin
        wt_pre_data_51 <= io_in_wt_data_51;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_52) begin
        wt_pre_data_52 <= io_in_wt_data_52;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_53) begin
        wt_pre_data_53 <= io_in_wt_data_53;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_54) begin
        wt_pre_data_54 <= io_in_wt_data_54;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_55) begin
        wt_pre_data_55 <= io_in_wt_data_55;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_56) begin
        wt_pre_data_56 <= io_in_wt_data_56;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_57) begin
        wt_pre_data_57 <= io_in_wt_data_57;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_58) begin
        wt_pre_data_58 <= io_in_wt_data_58;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_59) begin
        wt_pre_data_59 <= io_in_wt_data_59;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_60) begin
        wt_pre_data_60 <= io_in_wt_data_60;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_61) begin
        wt_pre_data_61 <= io_in_wt_data_61;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_62) begin
        wt_pre_data_62 <= io_in_wt_data_62;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_63) begin
        wt_pre_data_63 <= io_in_wt_data_63;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_64) begin
        wt_pre_data_64 <= io_in_wt_data_64;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_65) begin
        wt_pre_data_65 <= io_in_wt_data_65;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_66) begin
        wt_pre_data_66 <= io_in_wt_data_66;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_67) begin
        wt_pre_data_67 <= io_in_wt_data_67;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_68) begin
        wt_pre_data_68 <= io_in_wt_data_68;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_69) begin
        wt_pre_data_69 <= io_in_wt_data_69;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_70) begin
        wt_pre_data_70 <= io_in_wt_data_70;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_71) begin
        wt_pre_data_71 <= io_in_wt_data_71;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_72) begin
        wt_pre_data_72 <= io_in_wt_data_72;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_73) begin
        wt_pre_data_73 <= io_in_wt_data_73;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_74) begin
        wt_pre_data_74 <= io_in_wt_data_74;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_75) begin
        wt_pre_data_75 <= io_in_wt_data_75;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_76) begin
        wt_pre_data_76 <= io_in_wt_data_76;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_77) begin
        wt_pre_data_77 <= io_in_wt_data_77;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_78) begin
        wt_pre_data_78 <= io_in_wt_data_78;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_79) begin
        wt_pre_data_79 <= io_in_wt_data_79;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_80) begin
        wt_pre_data_80 <= io_in_wt_data_80;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_81) begin
        wt_pre_data_81 <= io_in_wt_data_81;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_82) begin
        wt_pre_data_82 <= io_in_wt_data_82;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_83) begin
        wt_pre_data_83 <= io_in_wt_data_83;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_84) begin
        wt_pre_data_84 <= io_in_wt_data_84;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_85) begin
        wt_pre_data_85 <= io_in_wt_data_85;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_86) begin
        wt_pre_data_86 <= io_in_wt_data_86;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_87) begin
        wt_pre_data_87 <= io_in_wt_data_87;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_88) begin
        wt_pre_data_88 <= io_in_wt_data_88;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_89) begin
        wt_pre_data_89 <= io_in_wt_data_89;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_90) begin
        wt_pre_data_90 <= io_in_wt_data_90;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_91) begin
        wt_pre_data_91 <= io_in_wt_data_91;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_92) begin
        wt_pre_data_92 <= io_in_wt_data_92;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_93) begin
        wt_pre_data_93 <= io_in_wt_data_93;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_94) begin
        wt_pre_data_94 <= io_in_wt_data_94;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_95) begin
        wt_pre_data_95 <= io_in_wt_data_95;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_96) begin
        wt_pre_data_96 <= io_in_wt_data_96;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_97) begin
        wt_pre_data_97 <= io_in_wt_data_97;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_98) begin
        wt_pre_data_98 <= io_in_wt_data_98;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_99) begin
        wt_pre_data_99 <= io_in_wt_data_99;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_100) begin
        wt_pre_data_100 <= io_in_wt_data_100;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_101) begin
        wt_pre_data_101 <= io_in_wt_data_101;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_102) begin
        wt_pre_data_102 <= io_in_wt_data_102;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_103) begin
        wt_pre_data_103 <= io_in_wt_data_103;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_104) begin
        wt_pre_data_104 <= io_in_wt_data_104;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_105) begin
        wt_pre_data_105 <= io_in_wt_data_105;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_106) begin
        wt_pre_data_106 <= io_in_wt_data_106;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_107) begin
        wt_pre_data_107 <= io_in_wt_data_107;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_108) begin
        wt_pre_data_108 <= io_in_wt_data_108;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_109) begin
        wt_pre_data_109 <= io_in_wt_data_109;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_110) begin
        wt_pre_data_110 <= io_in_wt_data_110;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_111) begin
        wt_pre_data_111 <= io_in_wt_data_111;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_112) begin
        wt_pre_data_112 <= io_in_wt_data_112;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_113) begin
        wt_pre_data_113 <= io_in_wt_data_113;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_114) begin
        wt_pre_data_114 <= io_in_wt_data_114;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_115) begin
        wt_pre_data_115 <= io_in_wt_data_115;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_116) begin
        wt_pre_data_116 <= io_in_wt_data_116;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_117) begin
        wt_pre_data_117 <= io_in_wt_data_117;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_118) begin
        wt_pre_data_118 <= io_in_wt_data_118;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_119) begin
        wt_pre_data_119 <= io_in_wt_data_119;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_120) begin
        wt_pre_data_120 <= io_in_wt_data_120;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_121) begin
        wt_pre_data_121 <= io_in_wt_data_121;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_122) begin
        wt_pre_data_122 <= io_in_wt_data_122;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_123) begin
        wt_pre_data_123 <= io_in_wt_data_123;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_124) begin
        wt_pre_data_124 <= io_in_wt_data_124;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_125) begin
        wt_pre_data_125 <= io_in_wt_data_125;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_126) begin
        wt_pre_data_126 <= io_in_wt_data_126;
      end
    end
    if (io_in_wt_pvld) begin
      if (io_in_wt_mask_127) begin
        wt_pre_data_127 <= io_in_wt_data_127;
      end
    end
    if (reset) begin
      wt_pre_sel_0 <= 1'h0;
    end else begin
      if (io_in_wt_pvld) begin
        wt_pre_sel_0 <= io_in_wt_sel_0;
      end
    end
    if (reset) begin
      dat_pre_nz_0 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_0 <= io_in_dat_mask_0;
      end
    end
    if (reset) begin
      dat_pre_nz_1 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_1 <= io_in_dat_mask_1;
      end
    end
    if (reset) begin
      dat_pre_nz_2 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_2 <= io_in_dat_mask_2;
      end
    end
    if (reset) begin
      dat_pre_nz_3 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_3 <= io_in_dat_mask_3;
      end
    end
    if (reset) begin
      dat_pre_nz_4 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_4 <= io_in_dat_mask_4;
      end
    end
    if (reset) begin
      dat_pre_nz_5 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_5 <= io_in_dat_mask_5;
      end
    end
    if (reset) begin
      dat_pre_nz_6 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_6 <= io_in_dat_mask_6;
      end
    end
    if (reset) begin
      dat_pre_nz_7 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_7 <= io_in_dat_mask_7;
      end
    end
    if (reset) begin
      dat_pre_nz_8 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_8 <= io_in_dat_mask_8;
      end
    end
    if (reset) begin
      dat_pre_nz_9 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_9 <= io_in_dat_mask_9;
      end
    end
    if (reset) begin
      dat_pre_nz_10 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_10 <= io_in_dat_mask_10;
      end
    end
    if (reset) begin
      dat_pre_nz_11 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_11 <= io_in_dat_mask_11;
      end
    end
    if (reset) begin
      dat_pre_nz_12 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_12 <= io_in_dat_mask_12;
      end
    end
    if (reset) begin
      dat_pre_nz_13 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_13 <= io_in_dat_mask_13;
      end
    end
    if (reset) begin
      dat_pre_nz_14 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_14 <= io_in_dat_mask_14;
      end
    end
    if (reset) begin
      dat_pre_nz_15 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_15 <= io_in_dat_mask_15;
      end
    end
    if (reset) begin
      dat_pre_nz_16 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_16 <= io_in_dat_mask_16;
      end
    end
    if (reset) begin
      dat_pre_nz_17 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_17 <= io_in_dat_mask_17;
      end
    end
    if (reset) begin
      dat_pre_nz_18 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_18 <= io_in_dat_mask_18;
      end
    end
    if (reset) begin
      dat_pre_nz_19 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_19 <= io_in_dat_mask_19;
      end
    end
    if (reset) begin
      dat_pre_nz_20 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_20 <= io_in_dat_mask_20;
      end
    end
    if (reset) begin
      dat_pre_nz_21 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_21 <= io_in_dat_mask_21;
      end
    end
    if (reset) begin
      dat_pre_nz_22 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_22 <= io_in_dat_mask_22;
      end
    end
    if (reset) begin
      dat_pre_nz_23 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_23 <= io_in_dat_mask_23;
      end
    end
    if (reset) begin
      dat_pre_nz_24 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_24 <= io_in_dat_mask_24;
      end
    end
    if (reset) begin
      dat_pre_nz_25 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_25 <= io_in_dat_mask_25;
      end
    end
    if (reset) begin
      dat_pre_nz_26 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_26 <= io_in_dat_mask_26;
      end
    end
    if (reset) begin
      dat_pre_nz_27 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_27 <= io_in_dat_mask_27;
      end
    end
    if (reset) begin
      dat_pre_nz_28 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_28 <= io_in_dat_mask_28;
      end
    end
    if (reset) begin
      dat_pre_nz_29 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_29 <= io_in_dat_mask_29;
      end
    end
    if (reset) begin
      dat_pre_nz_30 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_30 <= io_in_dat_mask_30;
      end
    end
    if (reset) begin
      dat_pre_nz_31 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_31 <= io_in_dat_mask_31;
      end
    end
    if (reset) begin
      dat_pre_nz_32 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_32 <= io_in_dat_mask_32;
      end
    end
    if (reset) begin
      dat_pre_nz_33 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_33 <= io_in_dat_mask_33;
      end
    end
    if (reset) begin
      dat_pre_nz_34 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_34 <= io_in_dat_mask_34;
      end
    end
    if (reset) begin
      dat_pre_nz_35 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_35 <= io_in_dat_mask_35;
      end
    end
    if (reset) begin
      dat_pre_nz_36 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_36 <= io_in_dat_mask_36;
      end
    end
    if (reset) begin
      dat_pre_nz_37 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_37 <= io_in_dat_mask_37;
      end
    end
    if (reset) begin
      dat_pre_nz_38 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_38 <= io_in_dat_mask_38;
      end
    end
    if (reset) begin
      dat_pre_nz_39 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_39 <= io_in_dat_mask_39;
      end
    end
    if (reset) begin
      dat_pre_nz_40 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_40 <= io_in_dat_mask_40;
      end
    end
    if (reset) begin
      dat_pre_nz_41 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_41 <= io_in_dat_mask_41;
      end
    end
    if (reset) begin
      dat_pre_nz_42 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_42 <= io_in_dat_mask_42;
      end
    end
    if (reset) begin
      dat_pre_nz_43 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_43 <= io_in_dat_mask_43;
      end
    end
    if (reset) begin
      dat_pre_nz_44 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_44 <= io_in_dat_mask_44;
      end
    end
    if (reset) begin
      dat_pre_nz_45 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_45 <= io_in_dat_mask_45;
      end
    end
    if (reset) begin
      dat_pre_nz_46 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_46 <= io_in_dat_mask_46;
      end
    end
    if (reset) begin
      dat_pre_nz_47 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_47 <= io_in_dat_mask_47;
      end
    end
    if (reset) begin
      dat_pre_nz_48 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_48 <= io_in_dat_mask_48;
      end
    end
    if (reset) begin
      dat_pre_nz_49 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_49 <= io_in_dat_mask_49;
      end
    end
    if (reset) begin
      dat_pre_nz_50 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_50 <= io_in_dat_mask_50;
      end
    end
    if (reset) begin
      dat_pre_nz_51 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_51 <= io_in_dat_mask_51;
      end
    end
    if (reset) begin
      dat_pre_nz_52 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_52 <= io_in_dat_mask_52;
      end
    end
    if (reset) begin
      dat_pre_nz_53 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_53 <= io_in_dat_mask_53;
      end
    end
    if (reset) begin
      dat_pre_nz_54 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_54 <= io_in_dat_mask_54;
      end
    end
    if (reset) begin
      dat_pre_nz_55 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_55 <= io_in_dat_mask_55;
      end
    end
    if (reset) begin
      dat_pre_nz_56 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_56 <= io_in_dat_mask_56;
      end
    end
    if (reset) begin
      dat_pre_nz_57 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_57 <= io_in_dat_mask_57;
      end
    end
    if (reset) begin
      dat_pre_nz_58 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_58 <= io_in_dat_mask_58;
      end
    end
    if (reset) begin
      dat_pre_nz_59 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_59 <= io_in_dat_mask_59;
      end
    end
    if (reset) begin
      dat_pre_nz_60 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_60 <= io_in_dat_mask_60;
      end
    end
    if (reset) begin
      dat_pre_nz_61 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_61 <= io_in_dat_mask_61;
      end
    end
    if (reset) begin
      dat_pre_nz_62 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_62 <= io_in_dat_mask_62;
      end
    end
    if (reset) begin
      dat_pre_nz_63 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_63 <= io_in_dat_mask_63;
      end
    end
    if (reset) begin
      dat_pre_nz_64 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_64 <= io_in_dat_mask_64;
      end
    end
    if (reset) begin
      dat_pre_nz_65 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_65 <= io_in_dat_mask_65;
      end
    end
    if (reset) begin
      dat_pre_nz_66 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_66 <= io_in_dat_mask_66;
      end
    end
    if (reset) begin
      dat_pre_nz_67 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_67 <= io_in_dat_mask_67;
      end
    end
    if (reset) begin
      dat_pre_nz_68 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_68 <= io_in_dat_mask_68;
      end
    end
    if (reset) begin
      dat_pre_nz_69 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_69 <= io_in_dat_mask_69;
      end
    end
    if (reset) begin
      dat_pre_nz_70 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_70 <= io_in_dat_mask_70;
      end
    end
    if (reset) begin
      dat_pre_nz_71 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_71 <= io_in_dat_mask_71;
      end
    end
    if (reset) begin
      dat_pre_nz_72 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_72 <= io_in_dat_mask_72;
      end
    end
    if (reset) begin
      dat_pre_nz_73 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_73 <= io_in_dat_mask_73;
      end
    end
    if (reset) begin
      dat_pre_nz_74 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_74 <= io_in_dat_mask_74;
      end
    end
    if (reset) begin
      dat_pre_nz_75 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_75 <= io_in_dat_mask_75;
      end
    end
    if (reset) begin
      dat_pre_nz_76 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_76 <= io_in_dat_mask_76;
      end
    end
    if (reset) begin
      dat_pre_nz_77 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_77 <= io_in_dat_mask_77;
      end
    end
    if (reset) begin
      dat_pre_nz_78 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_78 <= io_in_dat_mask_78;
      end
    end
    if (reset) begin
      dat_pre_nz_79 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_79 <= io_in_dat_mask_79;
      end
    end
    if (reset) begin
      dat_pre_nz_80 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_80 <= io_in_dat_mask_80;
      end
    end
    if (reset) begin
      dat_pre_nz_81 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_81 <= io_in_dat_mask_81;
      end
    end
    if (reset) begin
      dat_pre_nz_82 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_82 <= io_in_dat_mask_82;
      end
    end
    if (reset) begin
      dat_pre_nz_83 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_83 <= io_in_dat_mask_83;
      end
    end
    if (reset) begin
      dat_pre_nz_84 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_84 <= io_in_dat_mask_84;
      end
    end
    if (reset) begin
      dat_pre_nz_85 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_85 <= io_in_dat_mask_85;
      end
    end
    if (reset) begin
      dat_pre_nz_86 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_86 <= io_in_dat_mask_86;
      end
    end
    if (reset) begin
      dat_pre_nz_87 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_87 <= io_in_dat_mask_87;
      end
    end
    if (reset) begin
      dat_pre_nz_88 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_88 <= io_in_dat_mask_88;
      end
    end
    if (reset) begin
      dat_pre_nz_89 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_89 <= io_in_dat_mask_89;
      end
    end
    if (reset) begin
      dat_pre_nz_90 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_90 <= io_in_dat_mask_90;
      end
    end
    if (reset) begin
      dat_pre_nz_91 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_91 <= io_in_dat_mask_91;
      end
    end
    if (reset) begin
      dat_pre_nz_92 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_92 <= io_in_dat_mask_92;
      end
    end
    if (reset) begin
      dat_pre_nz_93 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_93 <= io_in_dat_mask_93;
      end
    end
    if (reset) begin
      dat_pre_nz_94 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_94 <= io_in_dat_mask_94;
      end
    end
    if (reset) begin
      dat_pre_nz_95 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_95 <= io_in_dat_mask_95;
      end
    end
    if (reset) begin
      dat_pre_nz_96 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_96 <= io_in_dat_mask_96;
      end
    end
    if (reset) begin
      dat_pre_nz_97 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_97 <= io_in_dat_mask_97;
      end
    end
    if (reset) begin
      dat_pre_nz_98 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_98 <= io_in_dat_mask_98;
      end
    end
    if (reset) begin
      dat_pre_nz_99 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_99 <= io_in_dat_mask_99;
      end
    end
    if (reset) begin
      dat_pre_nz_100 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_100 <= io_in_dat_mask_100;
      end
    end
    if (reset) begin
      dat_pre_nz_101 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_101 <= io_in_dat_mask_101;
      end
    end
    if (reset) begin
      dat_pre_nz_102 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_102 <= io_in_dat_mask_102;
      end
    end
    if (reset) begin
      dat_pre_nz_103 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_103 <= io_in_dat_mask_103;
      end
    end
    if (reset) begin
      dat_pre_nz_104 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_104 <= io_in_dat_mask_104;
      end
    end
    if (reset) begin
      dat_pre_nz_105 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_105 <= io_in_dat_mask_105;
      end
    end
    if (reset) begin
      dat_pre_nz_106 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_106 <= io_in_dat_mask_106;
      end
    end
    if (reset) begin
      dat_pre_nz_107 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_107 <= io_in_dat_mask_107;
      end
    end
    if (reset) begin
      dat_pre_nz_108 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_108 <= io_in_dat_mask_108;
      end
    end
    if (reset) begin
      dat_pre_nz_109 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_109 <= io_in_dat_mask_109;
      end
    end
    if (reset) begin
      dat_pre_nz_110 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_110 <= io_in_dat_mask_110;
      end
    end
    if (reset) begin
      dat_pre_nz_111 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_111 <= io_in_dat_mask_111;
      end
    end
    if (reset) begin
      dat_pre_nz_112 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_112 <= io_in_dat_mask_112;
      end
    end
    if (reset) begin
      dat_pre_nz_113 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_113 <= io_in_dat_mask_113;
      end
    end
    if (reset) begin
      dat_pre_nz_114 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_114 <= io_in_dat_mask_114;
      end
    end
    if (reset) begin
      dat_pre_nz_115 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_115 <= io_in_dat_mask_115;
      end
    end
    if (reset) begin
      dat_pre_nz_116 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_116 <= io_in_dat_mask_116;
      end
    end
    if (reset) begin
      dat_pre_nz_117 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_117 <= io_in_dat_mask_117;
      end
    end
    if (reset) begin
      dat_pre_nz_118 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_118 <= io_in_dat_mask_118;
      end
    end
    if (reset) begin
      dat_pre_nz_119 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_119 <= io_in_dat_mask_119;
      end
    end
    if (reset) begin
      dat_pre_nz_120 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_120 <= io_in_dat_mask_120;
      end
    end
    if (reset) begin
      dat_pre_nz_121 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_121 <= io_in_dat_mask_121;
      end
    end
    if (reset) begin
      dat_pre_nz_122 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_122 <= io_in_dat_mask_122;
      end
    end
    if (reset) begin
      dat_pre_nz_123 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_123 <= io_in_dat_mask_123;
      end
    end
    if (reset) begin
      dat_pre_nz_124 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_124 <= io_in_dat_mask_124;
      end
    end
    if (reset) begin
      dat_pre_nz_125 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_125 <= io_in_dat_mask_125;
      end
    end
    if (reset) begin
      dat_pre_nz_126 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_126 <= io_in_dat_mask_126;
      end
    end
    if (reset) begin
      dat_pre_nz_127 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_nz_127 <= io_in_dat_mask_127;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_0) begin
        dat_pre_data_0 <= io_in_dat_data_0;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_1) begin
        dat_pre_data_1 <= io_in_dat_data_1;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_2) begin
        dat_pre_data_2 <= io_in_dat_data_2;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_3) begin
        dat_pre_data_3 <= io_in_dat_data_3;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_4) begin
        dat_pre_data_4 <= io_in_dat_data_4;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_5) begin
        dat_pre_data_5 <= io_in_dat_data_5;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_6) begin
        dat_pre_data_6 <= io_in_dat_data_6;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_7) begin
        dat_pre_data_7 <= io_in_dat_data_7;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_8) begin
        dat_pre_data_8 <= io_in_dat_data_8;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_9) begin
        dat_pre_data_9 <= io_in_dat_data_9;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_10) begin
        dat_pre_data_10 <= io_in_dat_data_10;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_11) begin
        dat_pre_data_11 <= io_in_dat_data_11;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_12) begin
        dat_pre_data_12 <= io_in_dat_data_12;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_13) begin
        dat_pre_data_13 <= io_in_dat_data_13;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_14) begin
        dat_pre_data_14 <= io_in_dat_data_14;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_15) begin
        dat_pre_data_15 <= io_in_dat_data_15;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_16) begin
        dat_pre_data_16 <= io_in_dat_data_16;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_17) begin
        dat_pre_data_17 <= io_in_dat_data_17;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_18) begin
        dat_pre_data_18 <= io_in_dat_data_18;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_19) begin
        dat_pre_data_19 <= io_in_dat_data_19;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_20) begin
        dat_pre_data_20 <= io_in_dat_data_20;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_21) begin
        dat_pre_data_21 <= io_in_dat_data_21;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_22) begin
        dat_pre_data_22 <= io_in_dat_data_22;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_23) begin
        dat_pre_data_23 <= io_in_dat_data_23;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_24) begin
        dat_pre_data_24 <= io_in_dat_data_24;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_25) begin
        dat_pre_data_25 <= io_in_dat_data_25;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_26) begin
        dat_pre_data_26 <= io_in_dat_data_26;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_27) begin
        dat_pre_data_27 <= io_in_dat_data_27;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_28) begin
        dat_pre_data_28 <= io_in_dat_data_28;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_29) begin
        dat_pre_data_29 <= io_in_dat_data_29;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_30) begin
        dat_pre_data_30 <= io_in_dat_data_30;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_31) begin
        dat_pre_data_31 <= io_in_dat_data_31;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_32) begin
        dat_pre_data_32 <= io_in_dat_data_32;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_33) begin
        dat_pre_data_33 <= io_in_dat_data_33;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_34) begin
        dat_pre_data_34 <= io_in_dat_data_34;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_35) begin
        dat_pre_data_35 <= io_in_dat_data_35;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_36) begin
        dat_pre_data_36 <= io_in_dat_data_36;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_37) begin
        dat_pre_data_37 <= io_in_dat_data_37;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_38) begin
        dat_pre_data_38 <= io_in_dat_data_38;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_39) begin
        dat_pre_data_39 <= io_in_dat_data_39;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_40) begin
        dat_pre_data_40 <= io_in_dat_data_40;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_41) begin
        dat_pre_data_41 <= io_in_dat_data_41;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_42) begin
        dat_pre_data_42 <= io_in_dat_data_42;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_43) begin
        dat_pre_data_43 <= io_in_dat_data_43;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_44) begin
        dat_pre_data_44 <= io_in_dat_data_44;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_45) begin
        dat_pre_data_45 <= io_in_dat_data_45;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_46) begin
        dat_pre_data_46 <= io_in_dat_data_46;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_47) begin
        dat_pre_data_47 <= io_in_dat_data_47;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_48) begin
        dat_pre_data_48 <= io_in_dat_data_48;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_49) begin
        dat_pre_data_49 <= io_in_dat_data_49;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_50) begin
        dat_pre_data_50 <= io_in_dat_data_50;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_51) begin
        dat_pre_data_51 <= io_in_dat_data_51;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_52) begin
        dat_pre_data_52 <= io_in_dat_data_52;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_53) begin
        dat_pre_data_53 <= io_in_dat_data_53;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_54) begin
        dat_pre_data_54 <= io_in_dat_data_54;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_55) begin
        dat_pre_data_55 <= io_in_dat_data_55;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_56) begin
        dat_pre_data_56 <= io_in_dat_data_56;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_57) begin
        dat_pre_data_57 <= io_in_dat_data_57;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_58) begin
        dat_pre_data_58 <= io_in_dat_data_58;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_59) begin
        dat_pre_data_59 <= io_in_dat_data_59;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_60) begin
        dat_pre_data_60 <= io_in_dat_data_60;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_61) begin
        dat_pre_data_61 <= io_in_dat_data_61;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_62) begin
        dat_pre_data_62 <= io_in_dat_data_62;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_63) begin
        dat_pre_data_63 <= io_in_dat_data_63;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_64) begin
        dat_pre_data_64 <= io_in_dat_data_64;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_65) begin
        dat_pre_data_65 <= io_in_dat_data_65;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_66) begin
        dat_pre_data_66 <= io_in_dat_data_66;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_67) begin
        dat_pre_data_67 <= io_in_dat_data_67;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_68) begin
        dat_pre_data_68 <= io_in_dat_data_68;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_69) begin
        dat_pre_data_69 <= io_in_dat_data_69;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_70) begin
        dat_pre_data_70 <= io_in_dat_data_70;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_71) begin
        dat_pre_data_71 <= io_in_dat_data_71;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_72) begin
        dat_pre_data_72 <= io_in_dat_data_72;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_73) begin
        dat_pre_data_73 <= io_in_dat_data_73;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_74) begin
        dat_pre_data_74 <= io_in_dat_data_74;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_75) begin
        dat_pre_data_75 <= io_in_dat_data_75;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_76) begin
        dat_pre_data_76 <= io_in_dat_data_76;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_77) begin
        dat_pre_data_77 <= io_in_dat_data_77;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_78) begin
        dat_pre_data_78 <= io_in_dat_data_78;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_79) begin
        dat_pre_data_79 <= io_in_dat_data_79;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_80) begin
        dat_pre_data_80 <= io_in_dat_data_80;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_81) begin
        dat_pre_data_81 <= io_in_dat_data_81;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_82) begin
        dat_pre_data_82 <= io_in_dat_data_82;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_83) begin
        dat_pre_data_83 <= io_in_dat_data_83;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_84) begin
        dat_pre_data_84 <= io_in_dat_data_84;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_85) begin
        dat_pre_data_85 <= io_in_dat_data_85;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_86) begin
        dat_pre_data_86 <= io_in_dat_data_86;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_87) begin
        dat_pre_data_87 <= io_in_dat_data_87;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_88) begin
        dat_pre_data_88 <= io_in_dat_data_88;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_89) begin
        dat_pre_data_89 <= io_in_dat_data_89;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_90) begin
        dat_pre_data_90 <= io_in_dat_data_90;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_91) begin
        dat_pre_data_91 <= io_in_dat_data_91;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_92) begin
        dat_pre_data_92 <= io_in_dat_data_92;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_93) begin
        dat_pre_data_93 <= io_in_dat_data_93;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_94) begin
        dat_pre_data_94 <= io_in_dat_data_94;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_95) begin
        dat_pre_data_95 <= io_in_dat_data_95;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_96) begin
        dat_pre_data_96 <= io_in_dat_data_96;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_97) begin
        dat_pre_data_97 <= io_in_dat_data_97;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_98) begin
        dat_pre_data_98 <= io_in_dat_data_98;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_99) begin
        dat_pre_data_99 <= io_in_dat_data_99;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_100) begin
        dat_pre_data_100 <= io_in_dat_data_100;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_101) begin
        dat_pre_data_101 <= io_in_dat_data_101;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_102) begin
        dat_pre_data_102 <= io_in_dat_data_102;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_103) begin
        dat_pre_data_103 <= io_in_dat_data_103;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_104) begin
        dat_pre_data_104 <= io_in_dat_data_104;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_105) begin
        dat_pre_data_105 <= io_in_dat_data_105;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_106) begin
        dat_pre_data_106 <= io_in_dat_data_106;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_107) begin
        dat_pre_data_107 <= io_in_dat_data_107;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_108) begin
        dat_pre_data_108 <= io_in_dat_data_108;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_109) begin
        dat_pre_data_109 <= io_in_dat_data_109;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_110) begin
        dat_pre_data_110 <= io_in_dat_data_110;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_111) begin
        dat_pre_data_111 <= io_in_dat_data_111;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_112) begin
        dat_pre_data_112 <= io_in_dat_data_112;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_113) begin
        dat_pre_data_113 <= io_in_dat_data_113;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_114) begin
        dat_pre_data_114 <= io_in_dat_data_114;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_115) begin
        dat_pre_data_115 <= io_in_dat_data_115;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_116) begin
        dat_pre_data_116 <= io_in_dat_data_116;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_117) begin
        dat_pre_data_117 <= io_in_dat_data_117;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_118) begin
        dat_pre_data_118 <= io_in_dat_data_118;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_119) begin
        dat_pre_data_119 <= io_in_dat_data_119;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_120) begin
        dat_pre_data_120 <= io_in_dat_data_120;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_121) begin
        dat_pre_data_121 <= io_in_dat_data_121;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_122) begin
        dat_pre_data_122 <= io_in_dat_data_122;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_123) begin
        dat_pre_data_123 <= io_in_dat_data_123;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_124) begin
        dat_pre_data_124 <= io_in_dat_data_124;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_125) begin
        dat_pre_data_125 <= io_in_dat_data_125;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_126) begin
        dat_pre_data_126 <= io_in_dat_data_126;
      end
    end
    if (io_in_dat_pvld) begin
      if (io_in_dat_mask_127) begin
        dat_pre_data_127 <= io_in_dat_data_127;
      end
    end
    if (reset) begin
      dat_pre_pvld <= 1'h0;
    end else begin
      dat_pre_pvld <= io_in_dat_pvld;
    end
    if (reset) begin
      dat_pre_stripe_st_out_0 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_stripe_st_out_0 <= io_in_dat_stripe_st;
      end
    end
    if (reset) begin
      dat_pre_stripe_end_out_0 <= 1'h0;
    end else begin
      if (io_in_dat_pvld) begin
        dat_pre_stripe_end_out_0 <= io_in_dat_stripe_end;
      end
    end
    if (reset) begin
      wt_sd_pvld_0 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_pvld_0 <= 1'h1;
      end else begin
        if (dat_pre_stripe_st_out_0) begin
          wt_sd_pvld_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      wt_sd_nz_0_0 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_0 <= wt_pre_nz_0;
      end
    end
    if (reset) begin
      wt_sd_nz_0_1 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_1 <= wt_pre_nz_1;
      end
    end
    if (reset) begin
      wt_sd_nz_0_2 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_2 <= wt_pre_nz_2;
      end
    end
    if (reset) begin
      wt_sd_nz_0_3 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_3 <= wt_pre_nz_3;
      end
    end
    if (reset) begin
      wt_sd_nz_0_4 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_4 <= wt_pre_nz_4;
      end
    end
    if (reset) begin
      wt_sd_nz_0_5 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_5 <= wt_pre_nz_5;
      end
    end
    if (reset) begin
      wt_sd_nz_0_6 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_6 <= wt_pre_nz_6;
      end
    end
    if (reset) begin
      wt_sd_nz_0_7 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_7 <= wt_pre_nz_7;
      end
    end
    if (reset) begin
      wt_sd_nz_0_8 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_8 <= wt_pre_nz_8;
      end
    end
    if (reset) begin
      wt_sd_nz_0_9 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_9 <= wt_pre_nz_9;
      end
    end
    if (reset) begin
      wt_sd_nz_0_10 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_10 <= wt_pre_nz_10;
      end
    end
    if (reset) begin
      wt_sd_nz_0_11 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_11 <= wt_pre_nz_11;
      end
    end
    if (reset) begin
      wt_sd_nz_0_12 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_12 <= wt_pre_nz_12;
      end
    end
    if (reset) begin
      wt_sd_nz_0_13 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_13 <= wt_pre_nz_13;
      end
    end
    if (reset) begin
      wt_sd_nz_0_14 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_14 <= wt_pre_nz_14;
      end
    end
    if (reset) begin
      wt_sd_nz_0_15 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_15 <= wt_pre_nz_15;
      end
    end
    if (reset) begin
      wt_sd_nz_0_16 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_16 <= wt_pre_nz_16;
      end
    end
    if (reset) begin
      wt_sd_nz_0_17 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_17 <= wt_pre_nz_17;
      end
    end
    if (reset) begin
      wt_sd_nz_0_18 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_18 <= wt_pre_nz_18;
      end
    end
    if (reset) begin
      wt_sd_nz_0_19 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_19 <= wt_pre_nz_19;
      end
    end
    if (reset) begin
      wt_sd_nz_0_20 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_20 <= wt_pre_nz_20;
      end
    end
    if (reset) begin
      wt_sd_nz_0_21 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_21 <= wt_pre_nz_21;
      end
    end
    if (reset) begin
      wt_sd_nz_0_22 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_22 <= wt_pre_nz_22;
      end
    end
    if (reset) begin
      wt_sd_nz_0_23 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_23 <= wt_pre_nz_23;
      end
    end
    if (reset) begin
      wt_sd_nz_0_24 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_24 <= wt_pre_nz_24;
      end
    end
    if (reset) begin
      wt_sd_nz_0_25 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_25 <= wt_pre_nz_25;
      end
    end
    if (reset) begin
      wt_sd_nz_0_26 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_26 <= wt_pre_nz_26;
      end
    end
    if (reset) begin
      wt_sd_nz_0_27 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_27 <= wt_pre_nz_27;
      end
    end
    if (reset) begin
      wt_sd_nz_0_28 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_28 <= wt_pre_nz_28;
      end
    end
    if (reset) begin
      wt_sd_nz_0_29 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_29 <= wt_pre_nz_29;
      end
    end
    if (reset) begin
      wt_sd_nz_0_30 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_30 <= wt_pre_nz_30;
      end
    end
    if (reset) begin
      wt_sd_nz_0_31 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_31 <= wt_pre_nz_31;
      end
    end
    if (reset) begin
      wt_sd_nz_0_32 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_32 <= wt_pre_nz_32;
      end
    end
    if (reset) begin
      wt_sd_nz_0_33 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_33 <= wt_pre_nz_33;
      end
    end
    if (reset) begin
      wt_sd_nz_0_34 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_34 <= wt_pre_nz_34;
      end
    end
    if (reset) begin
      wt_sd_nz_0_35 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_35 <= wt_pre_nz_35;
      end
    end
    if (reset) begin
      wt_sd_nz_0_36 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_36 <= wt_pre_nz_36;
      end
    end
    if (reset) begin
      wt_sd_nz_0_37 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_37 <= wt_pre_nz_37;
      end
    end
    if (reset) begin
      wt_sd_nz_0_38 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_38 <= wt_pre_nz_38;
      end
    end
    if (reset) begin
      wt_sd_nz_0_39 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_39 <= wt_pre_nz_39;
      end
    end
    if (reset) begin
      wt_sd_nz_0_40 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_40 <= wt_pre_nz_40;
      end
    end
    if (reset) begin
      wt_sd_nz_0_41 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_41 <= wt_pre_nz_41;
      end
    end
    if (reset) begin
      wt_sd_nz_0_42 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_42 <= wt_pre_nz_42;
      end
    end
    if (reset) begin
      wt_sd_nz_0_43 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_43 <= wt_pre_nz_43;
      end
    end
    if (reset) begin
      wt_sd_nz_0_44 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_44 <= wt_pre_nz_44;
      end
    end
    if (reset) begin
      wt_sd_nz_0_45 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_45 <= wt_pre_nz_45;
      end
    end
    if (reset) begin
      wt_sd_nz_0_46 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_46 <= wt_pre_nz_46;
      end
    end
    if (reset) begin
      wt_sd_nz_0_47 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_47 <= wt_pre_nz_47;
      end
    end
    if (reset) begin
      wt_sd_nz_0_48 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_48 <= wt_pre_nz_48;
      end
    end
    if (reset) begin
      wt_sd_nz_0_49 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_49 <= wt_pre_nz_49;
      end
    end
    if (reset) begin
      wt_sd_nz_0_50 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_50 <= wt_pre_nz_50;
      end
    end
    if (reset) begin
      wt_sd_nz_0_51 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_51 <= wt_pre_nz_51;
      end
    end
    if (reset) begin
      wt_sd_nz_0_52 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_52 <= wt_pre_nz_52;
      end
    end
    if (reset) begin
      wt_sd_nz_0_53 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_53 <= wt_pre_nz_53;
      end
    end
    if (reset) begin
      wt_sd_nz_0_54 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_54 <= wt_pre_nz_54;
      end
    end
    if (reset) begin
      wt_sd_nz_0_55 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_55 <= wt_pre_nz_55;
      end
    end
    if (reset) begin
      wt_sd_nz_0_56 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_56 <= wt_pre_nz_56;
      end
    end
    if (reset) begin
      wt_sd_nz_0_57 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_57 <= wt_pre_nz_57;
      end
    end
    if (reset) begin
      wt_sd_nz_0_58 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_58 <= wt_pre_nz_58;
      end
    end
    if (reset) begin
      wt_sd_nz_0_59 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_59 <= wt_pre_nz_59;
      end
    end
    if (reset) begin
      wt_sd_nz_0_60 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_60 <= wt_pre_nz_60;
      end
    end
    if (reset) begin
      wt_sd_nz_0_61 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_61 <= wt_pre_nz_61;
      end
    end
    if (reset) begin
      wt_sd_nz_0_62 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_62 <= wt_pre_nz_62;
      end
    end
    if (reset) begin
      wt_sd_nz_0_63 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_63 <= wt_pre_nz_63;
      end
    end
    if (reset) begin
      wt_sd_nz_0_64 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_64 <= wt_pre_nz_64;
      end
    end
    if (reset) begin
      wt_sd_nz_0_65 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_65 <= wt_pre_nz_65;
      end
    end
    if (reset) begin
      wt_sd_nz_0_66 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_66 <= wt_pre_nz_66;
      end
    end
    if (reset) begin
      wt_sd_nz_0_67 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_67 <= wt_pre_nz_67;
      end
    end
    if (reset) begin
      wt_sd_nz_0_68 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_68 <= wt_pre_nz_68;
      end
    end
    if (reset) begin
      wt_sd_nz_0_69 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_69 <= wt_pre_nz_69;
      end
    end
    if (reset) begin
      wt_sd_nz_0_70 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_70 <= wt_pre_nz_70;
      end
    end
    if (reset) begin
      wt_sd_nz_0_71 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_71 <= wt_pre_nz_71;
      end
    end
    if (reset) begin
      wt_sd_nz_0_72 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_72 <= wt_pre_nz_72;
      end
    end
    if (reset) begin
      wt_sd_nz_0_73 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_73 <= wt_pre_nz_73;
      end
    end
    if (reset) begin
      wt_sd_nz_0_74 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_74 <= wt_pre_nz_74;
      end
    end
    if (reset) begin
      wt_sd_nz_0_75 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_75 <= wt_pre_nz_75;
      end
    end
    if (reset) begin
      wt_sd_nz_0_76 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_76 <= wt_pre_nz_76;
      end
    end
    if (reset) begin
      wt_sd_nz_0_77 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_77 <= wt_pre_nz_77;
      end
    end
    if (reset) begin
      wt_sd_nz_0_78 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_78 <= wt_pre_nz_78;
      end
    end
    if (reset) begin
      wt_sd_nz_0_79 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_79 <= wt_pre_nz_79;
      end
    end
    if (reset) begin
      wt_sd_nz_0_80 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_80 <= wt_pre_nz_80;
      end
    end
    if (reset) begin
      wt_sd_nz_0_81 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_81 <= wt_pre_nz_81;
      end
    end
    if (reset) begin
      wt_sd_nz_0_82 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_82 <= wt_pre_nz_82;
      end
    end
    if (reset) begin
      wt_sd_nz_0_83 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_83 <= wt_pre_nz_83;
      end
    end
    if (reset) begin
      wt_sd_nz_0_84 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_84 <= wt_pre_nz_84;
      end
    end
    if (reset) begin
      wt_sd_nz_0_85 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_85 <= wt_pre_nz_85;
      end
    end
    if (reset) begin
      wt_sd_nz_0_86 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_86 <= wt_pre_nz_86;
      end
    end
    if (reset) begin
      wt_sd_nz_0_87 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_87 <= wt_pre_nz_87;
      end
    end
    if (reset) begin
      wt_sd_nz_0_88 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_88 <= wt_pre_nz_88;
      end
    end
    if (reset) begin
      wt_sd_nz_0_89 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_89 <= wt_pre_nz_89;
      end
    end
    if (reset) begin
      wt_sd_nz_0_90 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_90 <= wt_pre_nz_90;
      end
    end
    if (reset) begin
      wt_sd_nz_0_91 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_91 <= wt_pre_nz_91;
      end
    end
    if (reset) begin
      wt_sd_nz_0_92 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_92 <= wt_pre_nz_92;
      end
    end
    if (reset) begin
      wt_sd_nz_0_93 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_93 <= wt_pre_nz_93;
      end
    end
    if (reset) begin
      wt_sd_nz_0_94 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_94 <= wt_pre_nz_94;
      end
    end
    if (reset) begin
      wt_sd_nz_0_95 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_95 <= wt_pre_nz_95;
      end
    end
    if (reset) begin
      wt_sd_nz_0_96 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_96 <= wt_pre_nz_96;
      end
    end
    if (reset) begin
      wt_sd_nz_0_97 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_97 <= wt_pre_nz_97;
      end
    end
    if (reset) begin
      wt_sd_nz_0_98 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_98 <= wt_pre_nz_98;
      end
    end
    if (reset) begin
      wt_sd_nz_0_99 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_99 <= wt_pre_nz_99;
      end
    end
    if (reset) begin
      wt_sd_nz_0_100 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_100 <= wt_pre_nz_100;
      end
    end
    if (reset) begin
      wt_sd_nz_0_101 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_101 <= wt_pre_nz_101;
      end
    end
    if (reset) begin
      wt_sd_nz_0_102 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_102 <= wt_pre_nz_102;
      end
    end
    if (reset) begin
      wt_sd_nz_0_103 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_103 <= wt_pre_nz_103;
      end
    end
    if (reset) begin
      wt_sd_nz_0_104 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_104 <= wt_pre_nz_104;
      end
    end
    if (reset) begin
      wt_sd_nz_0_105 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_105 <= wt_pre_nz_105;
      end
    end
    if (reset) begin
      wt_sd_nz_0_106 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_106 <= wt_pre_nz_106;
      end
    end
    if (reset) begin
      wt_sd_nz_0_107 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_107 <= wt_pre_nz_107;
      end
    end
    if (reset) begin
      wt_sd_nz_0_108 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_108 <= wt_pre_nz_108;
      end
    end
    if (reset) begin
      wt_sd_nz_0_109 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_109 <= wt_pre_nz_109;
      end
    end
    if (reset) begin
      wt_sd_nz_0_110 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_110 <= wt_pre_nz_110;
      end
    end
    if (reset) begin
      wt_sd_nz_0_111 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_111 <= wt_pre_nz_111;
      end
    end
    if (reset) begin
      wt_sd_nz_0_112 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_112 <= wt_pre_nz_112;
      end
    end
    if (reset) begin
      wt_sd_nz_0_113 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_113 <= wt_pre_nz_113;
      end
    end
    if (reset) begin
      wt_sd_nz_0_114 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_114 <= wt_pre_nz_114;
      end
    end
    if (reset) begin
      wt_sd_nz_0_115 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_115 <= wt_pre_nz_115;
      end
    end
    if (reset) begin
      wt_sd_nz_0_116 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_116 <= wt_pre_nz_116;
      end
    end
    if (reset) begin
      wt_sd_nz_0_117 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_117 <= wt_pre_nz_117;
      end
    end
    if (reset) begin
      wt_sd_nz_0_118 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_118 <= wt_pre_nz_118;
      end
    end
    if (reset) begin
      wt_sd_nz_0_119 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_119 <= wt_pre_nz_119;
      end
    end
    if (reset) begin
      wt_sd_nz_0_120 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_120 <= wt_pre_nz_120;
      end
    end
    if (reset) begin
      wt_sd_nz_0_121 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_121 <= wt_pre_nz_121;
      end
    end
    if (reset) begin
      wt_sd_nz_0_122 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_122 <= wt_pre_nz_122;
      end
    end
    if (reset) begin
      wt_sd_nz_0_123 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_123 <= wt_pre_nz_123;
      end
    end
    if (reset) begin
      wt_sd_nz_0_124 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_124 <= wt_pre_nz_124;
      end
    end
    if (reset) begin
      wt_sd_nz_0_125 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_125 <= wt_pre_nz_125;
      end
    end
    if (reset) begin
      wt_sd_nz_0_126 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_126 <= wt_pre_nz_126;
      end
    end
    if (reset) begin
      wt_sd_nz_0_127 <= 1'h0;
    end else begin
      if (wt_pre_sel_0) begin
        wt_sd_nz_0_127 <= wt_pre_nz_127;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_0) begin
        wt_sd_data_0_0 <= wt_pre_data_0;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_1) begin
        wt_sd_data_0_1 <= wt_pre_data_1;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_2) begin
        wt_sd_data_0_2 <= wt_pre_data_2;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_3) begin
        wt_sd_data_0_3 <= wt_pre_data_3;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_4) begin
        wt_sd_data_0_4 <= wt_pre_data_4;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_5) begin
        wt_sd_data_0_5 <= wt_pre_data_5;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_6) begin
        wt_sd_data_0_6 <= wt_pre_data_6;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_7) begin
        wt_sd_data_0_7 <= wt_pre_data_7;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_8) begin
        wt_sd_data_0_8 <= wt_pre_data_8;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_9) begin
        wt_sd_data_0_9 <= wt_pre_data_9;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_10) begin
        wt_sd_data_0_10 <= wt_pre_data_10;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_11) begin
        wt_sd_data_0_11 <= wt_pre_data_11;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_12) begin
        wt_sd_data_0_12 <= wt_pre_data_12;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_13) begin
        wt_sd_data_0_13 <= wt_pre_data_13;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_14) begin
        wt_sd_data_0_14 <= wt_pre_data_14;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_15) begin
        wt_sd_data_0_15 <= wt_pre_data_15;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_16) begin
        wt_sd_data_0_16 <= wt_pre_data_16;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_17) begin
        wt_sd_data_0_17 <= wt_pre_data_17;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_18) begin
        wt_sd_data_0_18 <= wt_pre_data_18;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_19) begin
        wt_sd_data_0_19 <= wt_pre_data_19;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_20) begin
        wt_sd_data_0_20 <= wt_pre_data_20;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_21) begin
        wt_sd_data_0_21 <= wt_pre_data_21;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_22) begin
        wt_sd_data_0_22 <= wt_pre_data_22;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_23) begin
        wt_sd_data_0_23 <= wt_pre_data_23;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_24) begin
        wt_sd_data_0_24 <= wt_pre_data_24;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_25) begin
        wt_sd_data_0_25 <= wt_pre_data_25;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_26) begin
        wt_sd_data_0_26 <= wt_pre_data_26;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_27) begin
        wt_sd_data_0_27 <= wt_pre_data_27;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_28) begin
        wt_sd_data_0_28 <= wt_pre_data_28;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_29) begin
        wt_sd_data_0_29 <= wt_pre_data_29;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_30) begin
        wt_sd_data_0_30 <= wt_pre_data_30;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_31) begin
        wt_sd_data_0_31 <= wt_pre_data_31;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_32) begin
        wt_sd_data_0_32 <= wt_pre_data_32;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_33) begin
        wt_sd_data_0_33 <= wt_pre_data_33;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_34) begin
        wt_sd_data_0_34 <= wt_pre_data_34;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_35) begin
        wt_sd_data_0_35 <= wt_pre_data_35;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_36) begin
        wt_sd_data_0_36 <= wt_pre_data_36;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_37) begin
        wt_sd_data_0_37 <= wt_pre_data_37;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_38) begin
        wt_sd_data_0_38 <= wt_pre_data_38;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_39) begin
        wt_sd_data_0_39 <= wt_pre_data_39;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_40) begin
        wt_sd_data_0_40 <= wt_pre_data_40;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_41) begin
        wt_sd_data_0_41 <= wt_pre_data_41;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_42) begin
        wt_sd_data_0_42 <= wt_pre_data_42;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_43) begin
        wt_sd_data_0_43 <= wt_pre_data_43;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_44) begin
        wt_sd_data_0_44 <= wt_pre_data_44;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_45) begin
        wt_sd_data_0_45 <= wt_pre_data_45;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_46) begin
        wt_sd_data_0_46 <= wt_pre_data_46;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_47) begin
        wt_sd_data_0_47 <= wt_pre_data_47;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_48) begin
        wt_sd_data_0_48 <= wt_pre_data_48;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_49) begin
        wt_sd_data_0_49 <= wt_pre_data_49;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_50) begin
        wt_sd_data_0_50 <= wt_pre_data_50;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_51) begin
        wt_sd_data_0_51 <= wt_pre_data_51;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_52) begin
        wt_sd_data_0_52 <= wt_pre_data_52;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_53) begin
        wt_sd_data_0_53 <= wt_pre_data_53;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_54) begin
        wt_sd_data_0_54 <= wt_pre_data_54;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_55) begin
        wt_sd_data_0_55 <= wt_pre_data_55;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_56) begin
        wt_sd_data_0_56 <= wt_pre_data_56;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_57) begin
        wt_sd_data_0_57 <= wt_pre_data_57;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_58) begin
        wt_sd_data_0_58 <= wt_pre_data_58;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_59) begin
        wt_sd_data_0_59 <= wt_pre_data_59;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_60) begin
        wt_sd_data_0_60 <= wt_pre_data_60;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_61) begin
        wt_sd_data_0_61 <= wt_pre_data_61;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_62) begin
        wt_sd_data_0_62 <= wt_pre_data_62;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_63) begin
        wt_sd_data_0_63 <= wt_pre_data_63;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_64) begin
        wt_sd_data_0_64 <= wt_pre_data_64;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_65) begin
        wt_sd_data_0_65 <= wt_pre_data_65;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_66) begin
        wt_sd_data_0_66 <= wt_pre_data_66;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_67) begin
        wt_sd_data_0_67 <= wt_pre_data_67;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_68) begin
        wt_sd_data_0_68 <= wt_pre_data_68;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_69) begin
        wt_sd_data_0_69 <= wt_pre_data_69;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_70) begin
        wt_sd_data_0_70 <= wt_pre_data_70;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_71) begin
        wt_sd_data_0_71 <= wt_pre_data_71;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_72) begin
        wt_sd_data_0_72 <= wt_pre_data_72;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_73) begin
        wt_sd_data_0_73 <= wt_pre_data_73;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_74) begin
        wt_sd_data_0_74 <= wt_pre_data_74;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_75) begin
        wt_sd_data_0_75 <= wt_pre_data_75;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_76) begin
        wt_sd_data_0_76 <= wt_pre_data_76;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_77) begin
        wt_sd_data_0_77 <= wt_pre_data_77;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_78) begin
        wt_sd_data_0_78 <= wt_pre_data_78;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_79) begin
        wt_sd_data_0_79 <= wt_pre_data_79;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_80) begin
        wt_sd_data_0_80 <= wt_pre_data_80;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_81) begin
        wt_sd_data_0_81 <= wt_pre_data_81;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_82) begin
        wt_sd_data_0_82 <= wt_pre_data_82;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_83) begin
        wt_sd_data_0_83 <= wt_pre_data_83;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_84) begin
        wt_sd_data_0_84 <= wt_pre_data_84;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_85) begin
        wt_sd_data_0_85 <= wt_pre_data_85;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_86) begin
        wt_sd_data_0_86 <= wt_pre_data_86;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_87) begin
        wt_sd_data_0_87 <= wt_pre_data_87;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_88) begin
        wt_sd_data_0_88 <= wt_pre_data_88;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_89) begin
        wt_sd_data_0_89 <= wt_pre_data_89;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_90) begin
        wt_sd_data_0_90 <= wt_pre_data_90;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_91) begin
        wt_sd_data_0_91 <= wt_pre_data_91;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_92) begin
        wt_sd_data_0_92 <= wt_pre_data_92;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_93) begin
        wt_sd_data_0_93 <= wt_pre_data_93;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_94) begin
        wt_sd_data_0_94 <= wt_pre_data_94;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_95) begin
        wt_sd_data_0_95 <= wt_pre_data_95;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_96) begin
        wt_sd_data_0_96 <= wt_pre_data_96;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_97) begin
        wt_sd_data_0_97 <= wt_pre_data_97;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_98) begin
        wt_sd_data_0_98 <= wt_pre_data_98;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_99) begin
        wt_sd_data_0_99 <= wt_pre_data_99;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_100) begin
        wt_sd_data_0_100 <= wt_pre_data_100;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_101) begin
        wt_sd_data_0_101 <= wt_pre_data_101;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_102) begin
        wt_sd_data_0_102 <= wt_pre_data_102;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_103) begin
        wt_sd_data_0_103 <= wt_pre_data_103;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_104) begin
        wt_sd_data_0_104 <= wt_pre_data_104;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_105) begin
        wt_sd_data_0_105 <= wt_pre_data_105;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_106) begin
        wt_sd_data_0_106 <= wt_pre_data_106;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_107) begin
        wt_sd_data_0_107 <= wt_pre_data_107;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_108) begin
        wt_sd_data_0_108 <= wt_pre_data_108;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_109) begin
        wt_sd_data_0_109 <= wt_pre_data_109;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_110) begin
        wt_sd_data_0_110 <= wt_pre_data_110;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_111) begin
        wt_sd_data_0_111 <= wt_pre_data_111;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_112) begin
        wt_sd_data_0_112 <= wt_pre_data_112;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_113) begin
        wt_sd_data_0_113 <= wt_pre_data_113;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_114) begin
        wt_sd_data_0_114 <= wt_pre_data_114;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_115) begin
        wt_sd_data_0_115 <= wt_pre_data_115;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_116) begin
        wt_sd_data_0_116 <= wt_pre_data_116;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_117) begin
        wt_sd_data_0_117 <= wt_pre_data_117;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_118) begin
        wt_sd_data_0_118 <= wt_pre_data_118;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_119) begin
        wt_sd_data_0_119 <= wt_pre_data_119;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_120) begin
        wt_sd_data_0_120 <= wt_pre_data_120;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_121) begin
        wt_sd_data_0_121 <= wt_pre_data_121;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_122) begin
        wt_sd_data_0_122 <= wt_pre_data_122;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_123) begin
        wt_sd_data_0_123 <= wt_pre_data_123;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_124) begin
        wt_sd_data_0_124 <= wt_pre_data_124;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_125) begin
        wt_sd_data_0_125 <= wt_pre_data_125;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_126) begin
        wt_sd_data_0_126 <= wt_pre_data_126;
      end
    end
    if (wt_pre_sel_0) begin
      if (wt_pre_nz_127) begin
        wt_sd_data_0_127 <= wt_pre_data_127;
      end
    end
    if (reset) begin
      dat_actv_stripe_end_0 <= 1'h0;
    end else begin
      dat_actv_stripe_end_0 <= dat_pre_stripe_end_out_0;
    end
    if (reset) begin
      wt_actv_vld_0 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_vld_0 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_vld_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_0 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_0 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_0 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_0 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_1 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_1 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_1 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_1 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_2 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_2 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_2 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_2 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_3 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_3 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_3 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_3 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_4 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_4 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_4 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_4 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_5 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_5 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_5 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_5 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_6 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_6 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_6 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_6 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_7 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_7 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_7 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_7 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_8 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_8 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_8 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_8 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_9 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_9 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_9 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_9 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_10 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_10 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_10 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_10 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_11 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_11 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_11 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_11 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_12 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_12 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_12 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_12 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_13 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_13 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_13 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_13 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_14 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_14 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_14 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_14 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_15 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_15 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_15 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_15 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_16 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_16 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_16 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_16 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_17 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_17 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_17 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_17 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_18 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_18 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_18 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_18 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_19 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_19 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_19 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_19 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_20 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_20 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_20 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_20 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_21 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_21 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_21 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_21 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_22 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_22 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_22 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_22 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_23 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_23 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_23 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_23 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_24 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_24 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_24 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_24 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_25 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_25 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_25 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_25 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_26 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_26 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_26 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_26 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_27 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_27 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_27 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_27 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_28 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_28 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_28 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_28 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_29 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_29 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_29 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_29 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_30 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_30 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_30 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_30 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_31 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_31 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_31 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_31 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_32 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_32 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_32 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_32 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_33 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_33 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_33 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_33 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_34 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_34 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_34 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_34 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_35 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_35 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_35 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_35 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_36 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_36 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_36 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_36 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_37 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_37 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_37 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_37 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_38 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_38 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_38 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_38 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_39 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_39 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_39 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_39 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_40 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_40 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_40 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_40 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_41 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_41 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_41 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_41 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_42 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_42 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_42 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_42 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_43 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_43 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_43 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_43 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_44 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_44 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_44 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_44 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_45 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_45 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_45 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_45 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_46 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_46 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_46 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_46 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_47 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_47 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_47 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_47 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_48 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_48 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_48 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_48 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_49 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_49 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_49 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_49 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_50 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_50 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_50 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_50 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_51 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_51 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_51 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_51 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_52 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_52 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_52 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_52 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_53 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_53 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_53 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_53 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_54 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_54 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_54 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_54 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_55 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_55 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_55 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_55 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_56 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_56 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_56 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_56 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_57 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_57 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_57 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_57 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_58 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_58 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_58 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_58 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_59 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_59 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_59 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_59 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_60 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_60 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_60 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_60 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_61 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_61 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_61 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_61 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_62 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_62 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_62 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_62 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_63 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_63 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_63 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_63 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_64 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_64 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_64 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_64 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_65 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_65 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_65 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_65 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_66 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_66 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_66 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_66 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_67 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_67 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_67 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_67 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_68 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_68 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_68 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_68 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_69 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_69 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_69 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_69 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_70 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_70 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_70 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_70 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_71 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_71 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_71 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_71 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_72 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_72 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_72 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_72 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_73 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_73 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_73 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_73 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_74 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_74 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_74 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_74 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_75 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_75 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_75 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_75 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_76 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_76 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_76 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_76 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_77 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_77 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_77 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_77 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_78 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_78 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_78 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_78 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_79 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_79 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_79 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_79 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_80 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_80 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_80 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_80 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_81 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_81 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_81 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_81 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_82 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_82 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_82 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_82 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_83 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_83 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_83 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_83 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_84 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_84 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_84 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_84 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_85 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_85 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_85 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_85 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_86 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_86 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_86 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_86 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_87 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_87 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_87 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_87 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_88 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_88 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_88 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_88 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_89 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_89 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_89 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_89 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_90 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_90 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_90 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_90 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_91 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_91 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_91 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_91 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_92 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_92 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_92 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_92 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_93 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_93 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_93 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_93 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_94 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_94 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_94 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_94 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_95 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_95 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_95 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_95 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_96 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_96 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_96 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_96 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_97 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_97 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_97 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_97 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_98 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_98 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_98 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_98 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_99 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_99 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_99 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_99 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_100 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_100 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_100 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_100 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_101 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_101 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_101 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_101 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_102 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_102 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_102 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_102 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_103 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_103 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_103 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_103 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_104 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_104 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_104 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_104 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_105 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_105 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_105 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_105 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_106 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_106 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_106 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_106 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_107 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_107 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_107 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_107 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_108 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_108 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_108 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_108 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_109 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_109 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_109 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_109 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_110 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_110 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_110 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_110 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_111 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_111 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_111 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_111 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_112 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_112 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_112 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_112 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_113 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_113 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_113 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_113 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_114 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_114 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_114 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_114 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_115 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_115 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_115 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_115 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_116 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_116 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_116 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_116 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_117 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_117 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_117 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_117 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_118 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_118 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_118 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_118 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_119 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_119 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_119 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_119 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_120 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_120 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_120 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_120 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_121 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_121 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_121 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_121 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_122 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_122 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_122 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_122 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_123 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_123 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_123 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_123 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_124 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_124 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_124 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_124 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_125 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_125 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_125 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_125 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_126 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_126 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_126 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_126 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_pvld_out_0_127 <= 1'h0;
    end else begin
      if (dat_pre_stripe_st_out_0) begin
        wt_actv_pvld_out_0_127 <= wt_sd_pvld_0;
      end else begin
        if (dat_actv_stripe_end_0) begin
          wt_actv_pvld_out_0_127 <= 1'h0;
        end else begin
          wt_actv_pvld_out_0_127 <= wt_actv_vld_0;
        end
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_0 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_0 <= wt_sd_nz_0_0;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_1 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_1 <= wt_sd_nz_0_1;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_2 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_2 <= wt_sd_nz_0_2;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_3 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_3 <= wt_sd_nz_0_3;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_4 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_4 <= wt_sd_nz_0_4;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_5 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_5 <= wt_sd_nz_0_5;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_6 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_6 <= wt_sd_nz_0_6;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_7 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_7 <= wt_sd_nz_0_7;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_8 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_8 <= wt_sd_nz_0_8;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_9 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_9 <= wt_sd_nz_0_9;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_10 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_10 <= wt_sd_nz_0_10;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_11 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_11 <= wt_sd_nz_0_11;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_12 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_12 <= wt_sd_nz_0_12;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_13 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_13 <= wt_sd_nz_0_13;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_14 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_14 <= wt_sd_nz_0_14;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_15 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_15 <= wt_sd_nz_0_15;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_16 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_16 <= wt_sd_nz_0_16;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_17 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_17 <= wt_sd_nz_0_17;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_18 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_18 <= wt_sd_nz_0_18;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_19 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_19 <= wt_sd_nz_0_19;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_20 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_20 <= wt_sd_nz_0_20;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_21 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_21 <= wt_sd_nz_0_21;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_22 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_22 <= wt_sd_nz_0_22;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_23 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_23 <= wt_sd_nz_0_23;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_24 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_24 <= wt_sd_nz_0_24;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_25 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_25 <= wt_sd_nz_0_25;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_26 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_26 <= wt_sd_nz_0_26;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_27 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_27 <= wt_sd_nz_0_27;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_28 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_28 <= wt_sd_nz_0_28;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_29 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_29 <= wt_sd_nz_0_29;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_30 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_30 <= wt_sd_nz_0_30;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_31 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_31 <= wt_sd_nz_0_31;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_32 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_32 <= wt_sd_nz_0_32;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_33 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_33 <= wt_sd_nz_0_33;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_34 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_34 <= wt_sd_nz_0_34;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_35 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_35 <= wt_sd_nz_0_35;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_36 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_36 <= wt_sd_nz_0_36;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_37 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_37 <= wt_sd_nz_0_37;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_38 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_38 <= wt_sd_nz_0_38;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_39 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_39 <= wt_sd_nz_0_39;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_40 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_40 <= wt_sd_nz_0_40;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_41 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_41 <= wt_sd_nz_0_41;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_42 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_42 <= wt_sd_nz_0_42;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_43 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_43 <= wt_sd_nz_0_43;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_44 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_44 <= wt_sd_nz_0_44;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_45 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_45 <= wt_sd_nz_0_45;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_46 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_46 <= wt_sd_nz_0_46;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_47 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_47 <= wt_sd_nz_0_47;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_48 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_48 <= wt_sd_nz_0_48;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_49 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_49 <= wt_sd_nz_0_49;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_50 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_50 <= wt_sd_nz_0_50;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_51 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_51 <= wt_sd_nz_0_51;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_52 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_52 <= wt_sd_nz_0_52;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_53 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_53 <= wt_sd_nz_0_53;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_54 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_54 <= wt_sd_nz_0_54;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_55 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_55 <= wt_sd_nz_0_55;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_56 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_56 <= wt_sd_nz_0_56;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_57 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_57 <= wt_sd_nz_0_57;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_58 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_58 <= wt_sd_nz_0_58;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_59 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_59 <= wt_sd_nz_0_59;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_60 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_60 <= wt_sd_nz_0_60;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_61 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_61 <= wt_sd_nz_0_61;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_62 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_62 <= wt_sd_nz_0_62;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_63 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_63 <= wt_sd_nz_0_63;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_64 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_64 <= wt_sd_nz_0_64;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_65 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_65 <= wt_sd_nz_0_65;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_66 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_66 <= wt_sd_nz_0_66;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_67 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_67 <= wt_sd_nz_0_67;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_68 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_68 <= wt_sd_nz_0_68;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_69 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_69 <= wt_sd_nz_0_69;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_70 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_70 <= wt_sd_nz_0_70;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_71 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_71 <= wt_sd_nz_0_71;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_72 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_72 <= wt_sd_nz_0_72;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_73 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_73 <= wt_sd_nz_0_73;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_74 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_74 <= wt_sd_nz_0_74;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_75 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_75 <= wt_sd_nz_0_75;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_76 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_76 <= wt_sd_nz_0_76;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_77 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_77 <= wt_sd_nz_0_77;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_78 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_78 <= wt_sd_nz_0_78;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_79 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_79 <= wt_sd_nz_0_79;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_80 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_80 <= wt_sd_nz_0_80;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_81 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_81 <= wt_sd_nz_0_81;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_82 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_82 <= wt_sd_nz_0_82;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_83 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_83 <= wt_sd_nz_0_83;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_84 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_84 <= wt_sd_nz_0_84;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_85 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_85 <= wt_sd_nz_0_85;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_86 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_86 <= wt_sd_nz_0_86;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_87 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_87 <= wt_sd_nz_0_87;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_88 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_88 <= wt_sd_nz_0_88;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_89 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_89 <= wt_sd_nz_0_89;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_90 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_90 <= wt_sd_nz_0_90;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_91 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_91 <= wt_sd_nz_0_91;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_92 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_92 <= wt_sd_nz_0_92;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_93 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_93 <= wt_sd_nz_0_93;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_94 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_94 <= wt_sd_nz_0_94;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_95 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_95 <= wt_sd_nz_0_95;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_96 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_96 <= wt_sd_nz_0_96;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_97 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_97 <= wt_sd_nz_0_97;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_98 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_98 <= wt_sd_nz_0_98;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_99 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_99 <= wt_sd_nz_0_99;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_100 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_100 <= wt_sd_nz_0_100;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_101 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_101 <= wt_sd_nz_0_101;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_102 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_102 <= wt_sd_nz_0_102;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_103 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_103 <= wt_sd_nz_0_103;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_104 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_104 <= wt_sd_nz_0_104;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_105 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_105 <= wt_sd_nz_0_105;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_106 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_106 <= wt_sd_nz_0_106;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_107 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_107 <= wt_sd_nz_0_107;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_108 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_108 <= wt_sd_nz_0_108;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_109 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_109 <= wt_sd_nz_0_109;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_110 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_110 <= wt_sd_nz_0_110;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_111 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_111 <= wt_sd_nz_0_111;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_112 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_112 <= wt_sd_nz_0_112;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_113 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_113 <= wt_sd_nz_0_113;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_114 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_114 <= wt_sd_nz_0_114;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_115 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_115 <= wt_sd_nz_0_115;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_116 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_116 <= wt_sd_nz_0_116;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_117 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_117 <= wt_sd_nz_0_117;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_118 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_118 <= wt_sd_nz_0_118;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_119 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_119 <= wt_sd_nz_0_119;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_120 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_120 <= wt_sd_nz_0_120;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_121 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_121 <= wt_sd_nz_0_121;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_122 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_122 <= wt_sd_nz_0_122;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_123 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_123 <= wt_sd_nz_0_123;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_124 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_124 <= wt_sd_nz_0_124;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_125 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_125 <= wt_sd_nz_0_125;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_126 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_126 <= wt_sd_nz_0_126;
      end
    end
    if (reset) begin
      wt_actv_nz_out_0_127 <= 1'h0;
    end else begin
      if (_T_50633) begin
        wt_actv_nz_out_0_127 <= wt_sd_nz_0_127;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_0) begin
        wt_actv_data_out_0_0 <= wt_sd_data_0_0;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_1) begin
        wt_actv_data_out_0_1 <= wt_sd_data_0_1;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_2) begin
        wt_actv_data_out_0_2 <= wt_sd_data_0_2;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_3) begin
        wt_actv_data_out_0_3 <= wt_sd_data_0_3;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_4) begin
        wt_actv_data_out_0_4 <= wt_sd_data_0_4;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_5) begin
        wt_actv_data_out_0_5 <= wt_sd_data_0_5;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_6) begin
        wt_actv_data_out_0_6 <= wt_sd_data_0_6;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_7) begin
        wt_actv_data_out_0_7 <= wt_sd_data_0_7;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_8) begin
        wt_actv_data_out_0_8 <= wt_sd_data_0_8;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_9) begin
        wt_actv_data_out_0_9 <= wt_sd_data_0_9;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_10) begin
        wt_actv_data_out_0_10 <= wt_sd_data_0_10;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_11) begin
        wt_actv_data_out_0_11 <= wt_sd_data_0_11;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_12) begin
        wt_actv_data_out_0_12 <= wt_sd_data_0_12;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_13) begin
        wt_actv_data_out_0_13 <= wt_sd_data_0_13;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_14) begin
        wt_actv_data_out_0_14 <= wt_sd_data_0_14;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_15) begin
        wt_actv_data_out_0_15 <= wt_sd_data_0_15;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_16) begin
        wt_actv_data_out_0_16 <= wt_sd_data_0_16;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_17) begin
        wt_actv_data_out_0_17 <= wt_sd_data_0_17;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_18) begin
        wt_actv_data_out_0_18 <= wt_sd_data_0_18;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_19) begin
        wt_actv_data_out_0_19 <= wt_sd_data_0_19;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_20) begin
        wt_actv_data_out_0_20 <= wt_sd_data_0_20;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_21) begin
        wt_actv_data_out_0_21 <= wt_sd_data_0_21;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_22) begin
        wt_actv_data_out_0_22 <= wt_sd_data_0_22;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_23) begin
        wt_actv_data_out_0_23 <= wt_sd_data_0_23;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_24) begin
        wt_actv_data_out_0_24 <= wt_sd_data_0_24;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_25) begin
        wt_actv_data_out_0_25 <= wt_sd_data_0_25;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_26) begin
        wt_actv_data_out_0_26 <= wt_sd_data_0_26;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_27) begin
        wt_actv_data_out_0_27 <= wt_sd_data_0_27;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_28) begin
        wt_actv_data_out_0_28 <= wt_sd_data_0_28;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_29) begin
        wt_actv_data_out_0_29 <= wt_sd_data_0_29;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_30) begin
        wt_actv_data_out_0_30 <= wt_sd_data_0_30;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_31) begin
        wt_actv_data_out_0_31 <= wt_sd_data_0_31;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_32) begin
        wt_actv_data_out_0_32 <= wt_sd_data_0_32;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_33) begin
        wt_actv_data_out_0_33 <= wt_sd_data_0_33;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_34) begin
        wt_actv_data_out_0_34 <= wt_sd_data_0_34;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_35) begin
        wt_actv_data_out_0_35 <= wt_sd_data_0_35;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_36) begin
        wt_actv_data_out_0_36 <= wt_sd_data_0_36;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_37) begin
        wt_actv_data_out_0_37 <= wt_sd_data_0_37;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_38) begin
        wt_actv_data_out_0_38 <= wt_sd_data_0_38;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_39) begin
        wt_actv_data_out_0_39 <= wt_sd_data_0_39;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_40) begin
        wt_actv_data_out_0_40 <= wt_sd_data_0_40;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_41) begin
        wt_actv_data_out_0_41 <= wt_sd_data_0_41;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_42) begin
        wt_actv_data_out_0_42 <= wt_sd_data_0_42;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_43) begin
        wt_actv_data_out_0_43 <= wt_sd_data_0_43;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_44) begin
        wt_actv_data_out_0_44 <= wt_sd_data_0_44;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_45) begin
        wt_actv_data_out_0_45 <= wt_sd_data_0_45;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_46) begin
        wt_actv_data_out_0_46 <= wt_sd_data_0_46;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_47) begin
        wt_actv_data_out_0_47 <= wt_sd_data_0_47;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_48) begin
        wt_actv_data_out_0_48 <= wt_sd_data_0_48;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_49) begin
        wt_actv_data_out_0_49 <= wt_sd_data_0_49;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_50) begin
        wt_actv_data_out_0_50 <= wt_sd_data_0_50;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_51) begin
        wt_actv_data_out_0_51 <= wt_sd_data_0_51;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_52) begin
        wt_actv_data_out_0_52 <= wt_sd_data_0_52;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_53) begin
        wt_actv_data_out_0_53 <= wt_sd_data_0_53;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_54) begin
        wt_actv_data_out_0_54 <= wt_sd_data_0_54;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_55) begin
        wt_actv_data_out_0_55 <= wt_sd_data_0_55;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_56) begin
        wt_actv_data_out_0_56 <= wt_sd_data_0_56;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_57) begin
        wt_actv_data_out_0_57 <= wt_sd_data_0_57;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_58) begin
        wt_actv_data_out_0_58 <= wt_sd_data_0_58;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_59) begin
        wt_actv_data_out_0_59 <= wt_sd_data_0_59;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_60) begin
        wt_actv_data_out_0_60 <= wt_sd_data_0_60;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_61) begin
        wt_actv_data_out_0_61 <= wt_sd_data_0_61;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_62) begin
        wt_actv_data_out_0_62 <= wt_sd_data_0_62;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_63) begin
        wt_actv_data_out_0_63 <= wt_sd_data_0_63;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_64) begin
        wt_actv_data_out_0_64 <= wt_sd_data_0_64;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_65) begin
        wt_actv_data_out_0_65 <= wt_sd_data_0_65;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_66) begin
        wt_actv_data_out_0_66 <= wt_sd_data_0_66;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_67) begin
        wt_actv_data_out_0_67 <= wt_sd_data_0_67;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_68) begin
        wt_actv_data_out_0_68 <= wt_sd_data_0_68;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_69) begin
        wt_actv_data_out_0_69 <= wt_sd_data_0_69;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_70) begin
        wt_actv_data_out_0_70 <= wt_sd_data_0_70;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_71) begin
        wt_actv_data_out_0_71 <= wt_sd_data_0_71;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_72) begin
        wt_actv_data_out_0_72 <= wt_sd_data_0_72;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_73) begin
        wt_actv_data_out_0_73 <= wt_sd_data_0_73;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_74) begin
        wt_actv_data_out_0_74 <= wt_sd_data_0_74;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_75) begin
        wt_actv_data_out_0_75 <= wt_sd_data_0_75;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_76) begin
        wt_actv_data_out_0_76 <= wt_sd_data_0_76;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_77) begin
        wt_actv_data_out_0_77 <= wt_sd_data_0_77;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_78) begin
        wt_actv_data_out_0_78 <= wt_sd_data_0_78;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_79) begin
        wt_actv_data_out_0_79 <= wt_sd_data_0_79;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_80) begin
        wt_actv_data_out_0_80 <= wt_sd_data_0_80;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_81) begin
        wt_actv_data_out_0_81 <= wt_sd_data_0_81;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_82) begin
        wt_actv_data_out_0_82 <= wt_sd_data_0_82;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_83) begin
        wt_actv_data_out_0_83 <= wt_sd_data_0_83;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_84) begin
        wt_actv_data_out_0_84 <= wt_sd_data_0_84;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_85) begin
        wt_actv_data_out_0_85 <= wt_sd_data_0_85;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_86) begin
        wt_actv_data_out_0_86 <= wt_sd_data_0_86;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_87) begin
        wt_actv_data_out_0_87 <= wt_sd_data_0_87;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_88) begin
        wt_actv_data_out_0_88 <= wt_sd_data_0_88;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_89) begin
        wt_actv_data_out_0_89 <= wt_sd_data_0_89;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_90) begin
        wt_actv_data_out_0_90 <= wt_sd_data_0_90;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_91) begin
        wt_actv_data_out_0_91 <= wt_sd_data_0_91;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_92) begin
        wt_actv_data_out_0_92 <= wt_sd_data_0_92;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_93) begin
        wt_actv_data_out_0_93 <= wt_sd_data_0_93;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_94) begin
        wt_actv_data_out_0_94 <= wt_sd_data_0_94;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_95) begin
        wt_actv_data_out_0_95 <= wt_sd_data_0_95;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_96) begin
        wt_actv_data_out_0_96 <= wt_sd_data_0_96;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_97) begin
        wt_actv_data_out_0_97 <= wt_sd_data_0_97;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_98) begin
        wt_actv_data_out_0_98 <= wt_sd_data_0_98;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_99) begin
        wt_actv_data_out_0_99 <= wt_sd_data_0_99;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_100) begin
        wt_actv_data_out_0_100 <= wt_sd_data_0_100;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_101) begin
        wt_actv_data_out_0_101 <= wt_sd_data_0_101;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_102) begin
        wt_actv_data_out_0_102 <= wt_sd_data_0_102;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_103) begin
        wt_actv_data_out_0_103 <= wt_sd_data_0_103;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_104) begin
        wt_actv_data_out_0_104 <= wt_sd_data_0_104;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_105) begin
        wt_actv_data_out_0_105 <= wt_sd_data_0_105;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_106) begin
        wt_actv_data_out_0_106 <= wt_sd_data_0_106;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_107) begin
        wt_actv_data_out_0_107 <= wt_sd_data_0_107;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_108) begin
        wt_actv_data_out_0_108 <= wt_sd_data_0_108;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_109) begin
        wt_actv_data_out_0_109 <= wt_sd_data_0_109;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_110) begin
        wt_actv_data_out_0_110 <= wt_sd_data_0_110;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_111) begin
        wt_actv_data_out_0_111 <= wt_sd_data_0_111;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_112) begin
        wt_actv_data_out_0_112 <= wt_sd_data_0_112;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_113) begin
        wt_actv_data_out_0_113 <= wt_sd_data_0_113;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_114) begin
        wt_actv_data_out_0_114 <= wt_sd_data_0_114;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_115) begin
        wt_actv_data_out_0_115 <= wt_sd_data_0_115;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_116) begin
        wt_actv_data_out_0_116 <= wt_sd_data_0_116;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_117) begin
        wt_actv_data_out_0_117 <= wt_sd_data_0_117;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_118) begin
        wt_actv_data_out_0_118 <= wt_sd_data_0_118;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_119) begin
        wt_actv_data_out_0_119 <= wt_sd_data_0_119;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_120) begin
        wt_actv_data_out_0_120 <= wt_sd_data_0_120;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_121) begin
        wt_actv_data_out_0_121 <= wt_sd_data_0_121;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_122) begin
        wt_actv_data_out_0_122 <= wt_sd_data_0_122;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_123) begin
        wt_actv_data_out_0_123 <= wt_sd_data_0_123;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_124) begin
        wt_actv_data_out_0_124 <= wt_sd_data_0_124;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_125) begin
        wt_actv_data_out_0_125 <= wt_sd_data_0_125;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_126) begin
        wt_actv_data_out_0_126 <= wt_sd_data_0_126;
      end
    end
    if (_T_50633) begin
      if (wt_sd_nz_0_127) begin
        wt_actv_data_out_0_127 <= wt_sd_data_0_127;
      end
    end
    if (_T_73569) begin
      dat_actv_data_reg_0_0 <= dat_pre_data_0;
    end
    if (_T_73570) begin
      dat_actv_data_reg_0_1 <= dat_pre_data_1;
    end
    if (_T_73571) begin
      dat_actv_data_reg_0_2 <= dat_pre_data_2;
    end
    if (_T_73572) begin
      dat_actv_data_reg_0_3 <= dat_pre_data_3;
    end
    if (_T_73573) begin
      dat_actv_data_reg_0_4 <= dat_pre_data_4;
    end
    if (_T_73574) begin
      dat_actv_data_reg_0_5 <= dat_pre_data_5;
    end
    if (_T_73575) begin
      dat_actv_data_reg_0_6 <= dat_pre_data_6;
    end
    if (_T_73576) begin
      dat_actv_data_reg_0_7 <= dat_pre_data_7;
    end
    if (_T_73577) begin
      dat_actv_data_reg_0_8 <= dat_pre_data_8;
    end
    if (_T_73578) begin
      dat_actv_data_reg_0_9 <= dat_pre_data_9;
    end
    if (_T_73579) begin
      dat_actv_data_reg_0_10 <= dat_pre_data_10;
    end
    if (_T_73580) begin
      dat_actv_data_reg_0_11 <= dat_pre_data_11;
    end
    if (_T_73581) begin
      dat_actv_data_reg_0_12 <= dat_pre_data_12;
    end
    if (_T_73582) begin
      dat_actv_data_reg_0_13 <= dat_pre_data_13;
    end
    if (_T_73583) begin
      dat_actv_data_reg_0_14 <= dat_pre_data_14;
    end
    if (_T_73584) begin
      dat_actv_data_reg_0_15 <= dat_pre_data_15;
    end
    if (_T_73585) begin
      dat_actv_data_reg_0_16 <= dat_pre_data_16;
    end
    if (_T_73586) begin
      dat_actv_data_reg_0_17 <= dat_pre_data_17;
    end
    if (_T_73587) begin
      dat_actv_data_reg_0_18 <= dat_pre_data_18;
    end
    if (_T_73588) begin
      dat_actv_data_reg_0_19 <= dat_pre_data_19;
    end
    if (_T_73589) begin
      dat_actv_data_reg_0_20 <= dat_pre_data_20;
    end
    if (_T_73590) begin
      dat_actv_data_reg_0_21 <= dat_pre_data_21;
    end
    if (_T_73591) begin
      dat_actv_data_reg_0_22 <= dat_pre_data_22;
    end
    if (_T_73592) begin
      dat_actv_data_reg_0_23 <= dat_pre_data_23;
    end
    if (_T_73593) begin
      dat_actv_data_reg_0_24 <= dat_pre_data_24;
    end
    if (_T_73594) begin
      dat_actv_data_reg_0_25 <= dat_pre_data_25;
    end
    if (_T_73595) begin
      dat_actv_data_reg_0_26 <= dat_pre_data_26;
    end
    if (_T_73596) begin
      dat_actv_data_reg_0_27 <= dat_pre_data_27;
    end
    if (_T_73597) begin
      dat_actv_data_reg_0_28 <= dat_pre_data_28;
    end
    if (_T_73598) begin
      dat_actv_data_reg_0_29 <= dat_pre_data_29;
    end
    if (_T_73599) begin
      dat_actv_data_reg_0_30 <= dat_pre_data_30;
    end
    if (_T_73600) begin
      dat_actv_data_reg_0_31 <= dat_pre_data_31;
    end
    if (_T_73601) begin
      dat_actv_data_reg_0_32 <= dat_pre_data_32;
    end
    if (_T_73602) begin
      dat_actv_data_reg_0_33 <= dat_pre_data_33;
    end
    if (_T_73603) begin
      dat_actv_data_reg_0_34 <= dat_pre_data_34;
    end
    if (_T_73604) begin
      dat_actv_data_reg_0_35 <= dat_pre_data_35;
    end
    if (_T_73605) begin
      dat_actv_data_reg_0_36 <= dat_pre_data_36;
    end
    if (_T_73606) begin
      dat_actv_data_reg_0_37 <= dat_pre_data_37;
    end
    if (_T_73607) begin
      dat_actv_data_reg_0_38 <= dat_pre_data_38;
    end
    if (_T_73608) begin
      dat_actv_data_reg_0_39 <= dat_pre_data_39;
    end
    if (_T_73609) begin
      dat_actv_data_reg_0_40 <= dat_pre_data_40;
    end
    if (_T_73610) begin
      dat_actv_data_reg_0_41 <= dat_pre_data_41;
    end
    if (_T_73611) begin
      dat_actv_data_reg_0_42 <= dat_pre_data_42;
    end
    if (_T_73612) begin
      dat_actv_data_reg_0_43 <= dat_pre_data_43;
    end
    if (_T_73613) begin
      dat_actv_data_reg_0_44 <= dat_pre_data_44;
    end
    if (_T_73614) begin
      dat_actv_data_reg_0_45 <= dat_pre_data_45;
    end
    if (_T_73615) begin
      dat_actv_data_reg_0_46 <= dat_pre_data_46;
    end
    if (_T_73616) begin
      dat_actv_data_reg_0_47 <= dat_pre_data_47;
    end
    if (_T_73617) begin
      dat_actv_data_reg_0_48 <= dat_pre_data_48;
    end
    if (_T_73618) begin
      dat_actv_data_reg_0_49 <= dat_pre_data_49;
    end
    if (_T_73619) begin
      dat_actv_data_reg_0_50 <= dat_pre_data_50;
    end
    if (_T_73620) begin
      dat_actv_data_reg_0_51 <= dat_pre_data_51;
    end
    if (_T_73621) begin
      dat_actv_data_reg_0_52 <= dat_pre_data_52;
    end
    if (_T_73622) begin
      dat_actv_data_reg_0_53 <= dat_pre_data_53;
    end
    if (_T_73623) begin
      dat_actv_data_reg_0_54 <= dat_pre_data_54;
    end
    if (_T_73624) begin
      dat_actv_data_reg_0_55 <= dat_pre_data_55;
    end
    if (_T_73625) begin
      dat_actv_data_reg_0_56 <= dat_pre_data_56;
    end
    if (_T_73626) begin
      dat_actv_data_reg_0_57 <= dat_pre_data_57;
    end
    if (_T_73627) begin
      dat_actv_data_reg_0_58 <= dat_pre_data_58;
    end
    if (_T_73628) begin
      dat_actv_data_reg_0_59 <= dat_pre_data_59;
    end
    if (_T_73629) begin
      dat_actv_data_reg_0_60 <= dat_pre_data_60;
    end
    if (_T_73630) begin
      dat_actv_data_reg_0_61 <= dat_pre_data_61;
    end
    if (_T_73631) begin
      dat_actv_data_reg_0_62 <= dat_pre_data_62;
    end
    if (_T_73632) begin
      dat_actv_data_reg_0_63 <= dat_pre_data_63;
    end
    if (_T_73633) begin
      dat_actv_data_reg_0_64 <= dat_pre_data_64;
    end
    if (_T_73634) begin
      dat_actv_data_reg_0_65 <= dat_pre_data_65;
    end
    if (_T_73635) begin
      dat_actv_data_reg_0_66 <= dat_pre_data_66;
    end
    if (_T_73636) begin
      dat_actv_data_reg_0_67 <= dat_pre_data_67;
    end
    if (_T_73637) begin
      dat_actv_data_reg_0_68 <= dat_pre_data_68;
    end
    if (_T_73638) begin
      dat_actv_data_reg_0_69 <= dat_pre_data_69;
    end
    if (_T_73639) begin
      dat_actv_data_reg_0_70 <= dat_pre_data_70;
    end
    if (_T_73640) begin
      dat_actv_data_reg_0_71 <= dat_pre_data_71;
    end
    if (_T_73641) begin
      dat_actv_data_reg_0_72 <= dat_pre_data_72;
    end
    if (_T_73642) begin
      dat_actv_data_reg_0_73 <= dat_pre_data_73;
    end
    if (_T_73643) begin
      dat_actv_data_reg_0_74 <= dat_pre_data_74;
    end
    if (_T_73644) begin
      dat_actv_data_reg_0_75 <= dat_pre_data_75;
    end
    if (_T_73645) begin
      dat_actv_data_reg_0_76 <= dat_pre_data_76;
    end
    if (_T_73646) begin
      dat_actv_data_reg_0_77 <= dat_pre_data_77;
    end
    if (_T_73647) begin
      dat_actv_data_reg_0_78 <= dat_pre_data_78;
    end
    if (_T_73648) begin
      dat_actv_data_reg_0_79 <= dat_pre_data_79;
    end
    if (_T_73649) begin
      dat_actv_data_reg_0_80 <= dat_pre_data_80;
    end
    if (_T_73650) begin
      dat_actv_data_reg_0_81 <= dat_pre_data_81;
    end
    if (_T_73651) begin
      dat_actv_data_reg_0_82 <= dat_pre_data_82;
    end
    if (_T_73652) begin
      dat_actv_data_reg_0_83 <= dat_pre_data_83;
    end
    if (_T_73653) begin
      dat_actv_data_reg_0_84 <= dat_pre_data_84;
    end
    if (_T_73654) begin
      dat_actv_data_reg_0_85 <= dat_pre_data_85;
    end
    if (_T_73655) begin
      dat_actv_data_reg_0_86 <= dat_pre_data_86;
    end
    if (_T_73656) begin
      dat_actv_data_reg_0_87 <= dat_pre_data_87;
    end
    if (_T_73657) begin
      dat_actv_data_reg_0_88 <= dat_pre_data_88;
    end
    if (_T_73658) begin
      dat_actv_data_reg_0_89 <= dat_pre_data_89;
    end
    if (_T_73659) begin
      dat_actv_data_reg_0_90 <= dat_pre_data_90;
    end
    if (_T_73660) begin
      dat_actv_data_reg_0_91 <= dat_pre_data_91;
    end
    if (_T_73661) begin
      dat_actv_data_reg_0_92 <= dat_pre_data_92;
    end
    if (_T_73662) begin
      dat_actv_data_reg_0_93 <= dat_pre_data_93;
    end
    if (_T_73663) begin
      dat_actv_data_reg_0_94 <= dat_pre_data_94;
    end
    if (_T_73664) begin
      dat_actv_data_reg_0_95 <= dat_pre_data_95;
    end
    if (_T_73665) begin
      dat_actv_data_reg_0_96 <= dat_pre_data_96;
    end
    if (_T_73666) begin
      dat_actv_data_reg_0_97 <= dat_pre_data_97;
    end
    if (_T_73667) begin
      dat_actv_data_reg_0_98 <= dat_pre_data_98;
    end
    if (_T_73668) begin
      dat_actv_data_reg_0_99 <= dat_pre_data_99;
    end
    if (_T_73669) begin
      dat_actv_data_reg_0_100 <= dat_pre_data_100;
    end
    if (_T_73670) begin
      dat_actv_data_reg_0_101 <= dat_pre_data_101;
    end
    if (_T_73671) begin
      dat_actv_data_reg_0_102 <= dat_pre_data_102;
    end
    if (_T_73672) begin
      dat_actv_data_reg_0_103 <= dat_pre_data_103;
    end
    if (_T_73673) begin
      dat_actv_data_reg_0_104 <= dat_pre_data_104;
    end
    if (_T_73674) begin
      dat_actv_data_reg_0_105 <= dat_pre_data_105;
    end
    if (_T_73675) begin
      dat_actv_data_reg_0_106 <= dat_pre_data_106;
    end
    if (_T_73676) begin
      dat_actv_data_reg_0_107 <= dat_pre_data_107;
    end
    if (_T_73677) begin
      dat_actv_data_reg_0_108 <= dat_pre_data_108;
    end
    if (_T_73678) begin
      dat_actv_data_reg_0_109 <= dat_pre_data_109;
    end
    if (_T_73679) begin
      dat_actv_data_reg_0_110 <= dat_pre_data_110;
    end
    if (_T_73680) begin
      dat_actv_data_reg_0_111 <= dat_pre_data_111;
    end
    if (_T_73681) begin
      dat_actv_data_reg_0_112 <= dat_pre_data_112;
    end
    if (_T_73682) begin
      dat_actv_data_reg_0_113 <= dat_pre_data_113;
    end
    if (_T_73683) begin
      dat_actv_data_reg_0_114 <= dat_pre_data_114;
    end
    if (_T_73684) begin
      dat_actv_data_reg_0_115 <= dat_pre_data_115;
    end
    if (_T_73685) begin
      dat_actv_data_reg_0_116 <= dat_pre_data_116;
    end
    if (_T_73686) begin
      dat_actv_data_reg_0_117 <= dat_pre_data_117;
    end
    if (_T_73687) begin
      dat_actv_data_reg_0_118 <= dat_pre_data_118;
    end
    if (_T_73688) begin
      dat_actv_data_reg_0_119 <= dat_pre_data_119;
    end
    if (_T_73689) begin
      dat_actv_data_reg_0_120 <= dat_pre_data_120;
    end
    if (_T_73690) begin
      dat_actv_data_reg_0_121 <= dat_pre_data_121;
    end
    if (_T_73691) begin
      dat_actv_data_reg_0_122 <= dat_pre_data_122;
    end
    if (_T_73692) begin
      dat_actv_data_reg_0_123 <= dat_pre_data_123;
    end
    if (_T_73693) begin
      dat_actv_data_reg_0_124 <= dat_pre_data_124;
    end
    if (_T_73694) begin
      dat_actv_data_reg_0_125 <= dat_pre_data_125;
    end
    if (_T_73695) begin
      dat_actv_data_reg_0_126 <= dat_pre_data_126;
    end
    if (_T_73696) begin
      dat_actv_data_reg_0_127 <= dat_pre_data_127;
    end
    if (reset) begin
      dat_actv_nz_reg_0_0 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_0 <= dat_pre_nz_0;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_1 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_1 <= dat_pre_nz_1;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_2 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_2 <= dat_pre_nz_2;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_3 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_3 <= dat_pre_nz_3;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_4 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_4 <= dat_pre_nz_4;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_5 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_5 <= dat_pre_nz_5;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_6 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_6 <= dat_pre_nz_6;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_7 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_7 <= dat_pre_nz_7;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_8 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_8 <= dat_pre_nz_8;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_9 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_9 <= dat_pre_nz_9;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_10 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_10 <= dat_pre_nz_10;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_11 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_11 <= dat_pre_nz_11;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_12 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_12 <= dat_pre_nz_12;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_13 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_13 <= dat_pre_nz_13;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_14 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_14 <= dat_pre_nz_14;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_15 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_15 <= dat_pre_nz_15;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_16 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_16 <= dat_pre_nz_16;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_17 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_17 <= dat_pre_nz_17;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_18 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_18 <= dat_pre_nz_18;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_19 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_19 <= dat_pre_nz_19;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_20 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_20 <= dat_pre_nz_20;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_21 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_21 <= dat_pre_nz_21;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_22 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_22 <= dat_pre_nz_22;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_23 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_23 <= dat_pre_nz_23;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_24 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_24 <= dat_pre_nz_24;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_25 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_25 <= dat_pre_nz_25;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_26 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_26 <= dat_pre_nz_26;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_27 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_27 <= dat_pre_nz_27;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_28 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_28 <= dat_pre_nz_28;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_29 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_29 <= dat_pre_nz_29;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_30 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_30 <= dat_pre_nz_30;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_31 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_31 <= dat_pre_nz_31;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_32 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_32 <= dat_pre_nz_32;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_33 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_33 <= dat_pre_nz_33;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_34 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_34 <= dat_pre_nz_34;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_35 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_35 <= dat_pre_nz_35;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_36 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_36 <= dat_pre_nz_36;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_37 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_37 <= dat_pre_nz_37;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_38 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_38 <= dat_pre_nz_38;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_39 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_39 <= dat_pre_nz_39;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_40 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_40 <= dat_pre_nz_40;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_41 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_41 <= dat_pre_nz_41;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_42 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_42 <= dat_pre_nz_42;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_43 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_43 <= dat_pre_nz_43;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_44 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_44 <= dat_pre_nz_44;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_45 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_45 <= dat_pre_nz_45;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_46 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_46 <= dat_pre_nz_46;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_47 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_47 <= dat_pre_nz_47;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_48 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_48 <= dat_pre_nz_48;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_49 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_49 <= dat_pre_nz_49;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_50 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_50 <= dat_pre_nz_50;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_51 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_51 <= dat_pre_nz_51;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_52 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_52 <= dat_pre_nz_52;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_53 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_53 <= dat_pre_nz_53;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_54 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_54 <= dat_pre_nz_54;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_55 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_55 <= dat_pre_nz_55;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_56 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_56 <= dat_pre_nz_56;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_57 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_57 <= dat_pre_nz_57;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_58 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_58 <= dat_pre_nz_58;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_59 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_59 <= dat_pre_nz_59;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_60 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_60 <= dat_pre_nz_60;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_61 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_61 <= dat_pre_nz_61;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_62 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_62 <= dat_pre_nz_62;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_63 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_63 <= dat_pre_nz_63;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_64 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_64 <= dat_pre_nz_64;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_65 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_65 <= dat_pre_nz_65;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_66 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_66 <= dat_pre_nz_66;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_67 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_67 <= dat_pre_nz_67;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_68 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_68 <= dat_pre_nz_68;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_69 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_69 <= dat_pre_nz_69;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_70 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_70 <= dat_pre_nz_70;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_71 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_71 <= dat_pre_nz_71;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_72 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_72 <= dat_pre_nz_72;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_73 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_73 <= dat_pre_nz_73;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_74 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_74 <= dat_pre_nz_74;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_75 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_75 <= dat_pre_nz_75;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_76 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_76 <= dat_pre_nz_76;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_77 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_77 <= dat_pre_nz_77;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_78 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_78 <= dat_pre_nz_78;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_79 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_79 <= dat_pre_nz_79;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_80 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_80 <= dat_pre_nz_80;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_81 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_81 <= dat_pre_nz_81;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_82 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_82 <= dat_pre_nz_82;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_83 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_83 <= dat_pre_nz_83;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_84 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_84 <= dat_pre_nz_84;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_85 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_85 <= dat_pre_nz_85;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_86 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_86 <= dat_pre_nz_86;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_87 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_87 <= dat_pre_nz_87;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_88 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_88 <= dat_pre_nz_88;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_89 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_89 <= dat_pre_nz_89;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_90 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_90 <= dat_pre_nz_90;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_91 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_91 <= dat_pre_nz_91;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_92 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_92 <= dat_pre_nz_92;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_93 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_93 <= dat_pre_nz_93;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_94 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_94 <= dat_pre_nz_94;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_95 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_95 <= dat_pre_nz_95;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_96 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_96 <= dat_pre_nz_96;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_97 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_97 <= dat_pre_nz_97;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_98 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_98 <= dat_pre_nz_98;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_99 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_99 <= dat_pre_nz_99;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_100 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_100 <= dat_pre_nz_100;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_101 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_101 <= dat_pre_nz_101;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_102 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_102 <= dat_pre_nz_102;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_103 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_103 <= dat_pre_nz_103;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_104 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_104 <= dat_pre_nz_104;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_105 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_105 <= dat_pre_nz_105;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_106 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_106 <= dat_pre_nz_106;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_107 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_107 <= dat_pre_nz_107;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_108 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_108 <= dat_pre_nz_108;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_109 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_109 <= dat_pre_nz_109;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_110 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_110 <= dat_pre_nz_110;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_111 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_111 <= dat_pre_nz_111;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_112 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_112 <= dat_pre_nz_112;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_113 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_113 <= dat_pre_nz_113;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_114 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_114 <= dat_pre_nz_114;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_115 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_115 <= dat_pre_nz_115;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_116 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_116 <= dat_pre_nz_116;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_117 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_117 <= dat_pre_nz_117;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_118 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_118 <= dat_pre_nz_118;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_119 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_119 <= dat_pre_nz_119;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_120 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_120 <= dat_pre_nz_120;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_121 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_121 <= dat_pre_nz_121;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_122 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_122 <= dat_pre_nz_122;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_123 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_123 <= dat_pre_nz_123;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_124 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_124 <= dat_pre_nz_124;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_125 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_125 <= dat_pre_nz_125;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_126 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_126 <= dat_pre_nz_126;
      end
    end
    if (reset) begin
      dat_actv_nz_reg_0_127 <= 1'h0;
    end else begin
      if (dat_pre_pvld) begin
        dat_actv_nz_reg_0_127 <= dat_pre_nz_127;
      end
    end
    if (reset) begin
      dat_actv_pvld_reg_0_0 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_0 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_1 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_1 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_2 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_2 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_3 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_3 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_4 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_4 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_5 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_5 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_6 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_6 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_7 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_7 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_8 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_8 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_9 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_9 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_10 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_10 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_11 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_11 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_12 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_12 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_13 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_13 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_14 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_14 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_15 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_15 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_16 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_16 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_17 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_17 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_18 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_18 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_19 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_19 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_20 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_20 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_21 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_21 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_22 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_22 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_23 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_23 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_24 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_24 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_25 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_25 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_26 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_26 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_27 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_27 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_28 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_28 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_29 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_29 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_30 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_30 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_31 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_31 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_32 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_32 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_33 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_33 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_34 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_34 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_35 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_35 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_36 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_36 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_37 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_37 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_38 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_38 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_39 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_39 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_40 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_40 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_41 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_41 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_42 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_42 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_43 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_43 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_44 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_44 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_45 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_45 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_46 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_46 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_47 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_47 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_48 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_48 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_49 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_49 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_50 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_50 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_51 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_51 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_52 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_52 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_53 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_53 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_54 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_54 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_55 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_55 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_56 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_56 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_57 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_57 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_58 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_58 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_59 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_59 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_60 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_60 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_61 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_61 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_62 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_62 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_63 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_63 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_64 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_64 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_65 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_65 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_66 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_66 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_67 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_67 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_68 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_68 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_69 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_69 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_70 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_70 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_71 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_71 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_72 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_72 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_73 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_73 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_74 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_74 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_75 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_75 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_76 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_76 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_77 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_77 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_78 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_78 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_79 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_79 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_80 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_80 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_81 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_81 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_82 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_82 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_83 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_83 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_84 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_84 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_85 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_85 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_86 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_86 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_87 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_87 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_88 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_88 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_89 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_89 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_90 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_90 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_91 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_91 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_92 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_92 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_93 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_93 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_94 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_94 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_95 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_95 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_96 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_96 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_97 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_97 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_98 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_98 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_99 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_99 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_100 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_100 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_101 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_101 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_102 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_102 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_103 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_103 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_104 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_104 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_105 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_105 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_106 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_106 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_107 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_107 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_108 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_108 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_109 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_109 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_110 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_110 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_111 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_111 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_112 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_112 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_113 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_113 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_114 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_114 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_115 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_115 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_116 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_116 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_117 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_117 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_118 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_118 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_119 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_119 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_120 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_120 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_121 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_121 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_122 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_122 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_123 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_123 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_124 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_124 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_125 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_125 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_126 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_126 <= dat_pre_pvld;
    end
    if (reset) begin
      dat_actv_pvld_reg_0_127 <= 1'h0;
    end else begin
      dat_actv_pvld_reg_0_127 <= dat_pre_pvld;
    end
  end
endmodule
module NV_NVDLA_CMAC_CORE_mac(
  input         clock,
  input  [7:0]  io_dat_actv_data_0,
  input  [7:0]  io_dat_actv_data_1,
  input  [7:0]  io_dat_actv_data_2,
  input  [7:0]  io_dat_actv_data_3,
  input  [7:0]  io_dat_actv_data_4,
  input  [7:0]  io_dat_actv_data_5,
  input  [7:0]  io_dat_actv_data_6,
  input  [7:0]  io_dat_actv_data_7,
  input  [7:0]  io_dat_actv_data_8,
  input  [7:0]  io_dat_actv_data_9,
  input  [7:0]  io_dat_actv_data_10,
  input  [7:0]  io_dat_actv_data_11,
  input  [7:0]  io_dat_actv_data_12,
  input  [7:0]  io_dat_actv_data_13,
  input  [7:0]  io_dat_actv_data_14,
  input  [7:0]  io_dat_actv_data_15,
  input  [7:0]  io_dat_actv_data_16,
  input  [7:0]  io_dat_actv_data_17,
  input  [7:0]  io_dat_actv_data_18,
  input  [7:0]  io_dat_actv_data_19,
  input  [7:0]  io_dat_actv_data_20,
  input  [7:0]  io_dat_actv_data_21,
  input  [7:0]  io_dat_actv_data_22,
  input  [7:0]  io_dat_actv_data_23,
  input  [7:0]  io_dat_actv_data_24,
  input  [7:0]  io_dat_actv_data_25,
  input  [7:0]  io_dat_actv_data_26,
  input  [7:0]  io_dat_actv_data_27,
  input  [7:0]  io_dat_actv_data_28,
  input  [7:0]  io_dat_actv_data_29,
  input  [7:0]  io_dat_actv_data_30,
  input  [7:0]  io_dat_actv_data_31,
  input  [7:0]  io_dat_actv_data_32,
  input  [7:0]  io_dat_actv_data_33,
  input  [7:0]  io_dat_actv_data_34,
  input  [7:0]  io_dat_actv_data_35,
  input  [7:0]  io_dat_actv_data_36,
  input  [7:0]  io_dat_actv_data_37,
  input  [7:0]  io_dat_actv_data_38,
  input  [7:0]  io_dat_actv_data_39,
  input  [7:0]  io_dat_actv_data_40,
  input  [7:0]  io_dat_actv_data_41,
  input  [7:0]  io_dat_actv_data_42,
  input  [7:0]  io_dat_actv_data_43,
  input  [7:0]  io_dat_actv_data_44,
  input  [7:0]  io_dat_actv_data_45,
  input  [7:0]  io_dat_actv_data_46,
  input  [7:0]  io_dat_actv_data_47,
  input  [7:0]  io_dat_actv_data_48,
  input  [7:0]  io_dat_actv_data_49,
  input  [7:0]  io_dat_actv_data_50,
  input  [7:0]  io_dat_actv_data_51,
  input  [7:0]  io_dat_actv_data_52,
  input  [7:0]  io_dat_actv_data_53,
  input  [7:0]  io_dat_actv_data_54,
  input  [7:0]  io_dat_actv_data_55,
  input  [7:0]  io_dat_actv_data_56,
  input  [7:0]  io_dat_actv_data_57,
  input  [7:0]  io_dat_actv_data_58,
  input  [7:0]  io_dat_actv_data_59,
  input  [7:0]  io_dat_actv_data_60,
  input  [7:0]  io_dat_actv_data_61,
  input  [7:0]  io_dat_actv_data_62,
  input  [7:0]  io_dat_actv_data_63,
  input  [7:0]  io_dat_actv_data_64,
  input  [7:0]  io_dat_actv_data_65,
  input  [7:0]  io_dat_actv_data_66,
  input  [7:0]  io_dat_actv_data_67,
  input  [7:0]  io_dat_actv_data_68,
  input  [7:0]  io_dat_actv_data_69,
  input  [7:0]  io_dat_actv_data_70,
  input  [7:0]  io_dat_actv_data_71,
  input  [7:0]  io_dat_actv_data_72,
  input  [7:0]  io_dat_actv_data_73,
  input  [7:0]  io_dat_actv_data_74,
  input  [7:0]  io_dat_actv_data_75,
  input  [7:0]  io_dat_actv_data_76,
  input  [7:0]  io_dat_actv_data_77,
  input  [7:0]  io_dat_actv_data_78,
  input  [7:0]  io_dat_actv_data_79,
  input  [7:0]  io_dat_actv_data_80,
  input  [7:0]  io_dat_actv_data_81,
  input  [7:0]  io_dat_actv_data_82,
  input  [7:0]  io_dat_actv_data_83,
  input  [7:0]  io_dat_actv_data_84,
  input  [7:0]  io_dat_actv_data_85,
  input  [7:0]  io_dat_actv_data_86,
  input  [7:0]  io_dat_actv_data_87,
  input  [7:0]  io_dat_actv_data_88,
  input  [7:0]  io_dat_actv_data_89,
  input  [7:0]  io_dat_actv_data_90,
  input  [7:0]  io_dat_actv_data_91,
  input  [7:0]  io_dat_actv_data_92,
  input  [7:0]  io_dat_actv_data_93,
  input  [7:0]  io_dat_actv_data_94,
  input  [7:0]  io_dat_actv_data_95,
  input  [7:0]  io_dat_actv_data_96,
  input  [7:0]  io_dat_actv_data_97,
  input  [7:0]  io_dat_actv_data_98,
  input  [7:0]  io_dat_actv_data_99,
  input  [7:0]  io_dat_actv_data_100,
  input  [7:0]  io_dat_actv_data_101,
  input  [7:0]  io_dat_actv_data_102,
  input  [7:0]  io_dat_actv_data_103,
  input  [7:0]  io_dat_actv_data_104,
  input  [7:0]  io_dat_actv_data_105,
  input  [7:0]  io_dat_actv_data_106,
  input  [7:0]  io_dat_actv_data_107,
  input  [7:0]  io_dat_actv_data_108,
  input  [7:0]  io_dat_actv_data_109,
  input  [7:0]  io_dat_actv_data_110,
  input  [7:0]  io_dat_actv_data_111,
  input  [7:0]  io_dat_actv_data_112,
  input  [7:0]  io_dat_actv_data_113,
  input  [7:0]  io_dat_actv_data_114,
  input  [7:0]  io_dat_actv_data_115,
  input  [7:0]  io_dat_actv_data_116,
  input  [7:0]  io_dat_actv_data_117,
  input  [7:0]  io_dat_actv_data_118,
  input  [7:0]  io_dat_actv_data_119,
  input  [7:0]  io_dat_actv_data_120,
  input  [7:0]  io_dat_actv_data_121,
  input  [7:0]  io_dat_actv_data_122,
  input  [7:0]  io_dat_actv_data_123,
  input  [7:0]  io_dat_actv_data_124,
  input  [7:0]  io_dat_actv_data_125,
  input  [7:0]  io_dat_actv_data_126,
  input  [7:0]  io_dat_actv_data_127,
  input         io_dat_actv_nz_0,
  input         io_dat_actv_nz_1,
  input         io_dat_actv_nz_2,
  input         io_dat_actv_nz_3,
  input         io_dat_actv_nz_4,
  input         io_dat_actv_nz_5,
  input         io_dat_actv_nz_6,
  input         io_dat_actv_nz_7,
  input         io_dat_actv_nz_8,
  input         io_dat_actv_nz_9,
  input         io_dat_actv_nz_10,
  input         io_dat_actv_nz_11,
  input         io_dat_actv_nz_12,
  input         io_dat_actv_nz_13,
  input         io_dat_actv_nz_14,
  input         io_dat_actv_nz_15,
  input         io_dat_actv_nz_16,
  input         io_dat_actv_nz_17,
  input         io_dat_actv_nz_18,
  input         io_dat_actv_nz_19,
  input         io_dat_actv_nz_20,
  input         io_dat_actv_nz_21,
  input         io_dat_actv_nz_22,
  input         io_dat_actv_nz_23,
  input         io_dat_actv_nz_24,
  input         io_dat_actv_nz_25,
  input         io_dat_actv_nz_26,
  input         io_dat_actv_nz_27,
  input         io_dat_actv_nz_28,
  input         io_dat_actv_nz_29,
  input         io_dat_actv_nz_30,
  input         io_dat_actv_nz_31,
  input         io_dat_actv_nz_32,
  input         io_dat_actv_nz_33,
  input         io_dat_actv_nz_34,
  input         io_dat_actv_nz_35,
  input         io_dat_actv_nz_36,
  input         io_dat_actv_nz_37,
  input         io_dat_actv_nz_38,
  input         io_dat_actv_nz_39,
  input         io_dat_actv_nz_40,
  input         io_dat_actv_nz_41,
  input         io_dat_actv_nz_42,
  input         io_dat_actv_nz_43,
  input         io_dat_actv_nz_44,
  input         io_dat_actv_nz_45,
  input         io_dat_actv_nz_46,
  input         io_dat_actv_nz_47,
  input         io_dat_actv_nz_48,
  input         io_dat_actv_nz_49,
  input         io_dat_actv_nz_50,
  input         io_dat_actv_nz_51,
  input         io_dat_actv_nz_52,
  input         io_dat_actv_nz_53,
  input         io_dat_actv_nz_54,
  input         io_dat_actv_nz_55,
  input         io_dat_actv_nz_56,
  input         io_dat_actv_nz_57,
  input         io_dat_actv_nz_58,
  input         io_dat_actv_nz_59,
  input         io_dat_actv_nz_60,
  input         io_dat_actv_nz_61,
  input         io_dat_actv_nz_62,
  input         io_dat_actv_nz_63,
  input         io_dat_actv_nz_64,
  input         io_dat_actv_nz_65,
  input         io_dat_actv_nz_66,
  input         io_dat_actv_nz_67,
  input         io_dat_actv_nz_68,
  input         io_dat_actv_nz_69,
  input         io_dat_actv_nz_70,
  input         io_dat_actv_nz_71,
  input         io_dat_actv_nz_72,
  input         io_dat_actv_nz_73,
  input         io_dat_actv_nz_74,
  input         io_dat_actv_nz_75,
  input         io_dat_actv_nz_76,
  input         io_dat_actv_nz_77,
  input         io_dat_actv_nz_78,
  input         io_dat_actv_nz_79,
  input         io_dat_actv_nz_80,
  input         io_dat_actv_nz_81,
  input         io_dat_actv_nz_82,
  input         io_dat_actv_nz_83,
  input         io_dat_actv_nz_84,
  input         io_dat_actv_nz_85,
  input         io_dat_actv_nz_86,
  input         io_dat_actv_nz_87,
  input         io_dat_actv_nz_88,
  input         io_dat_actv_nz_89,
  input         io_dat_actv_nz_90,
  input         io_dat_actv_nz_91,
  input         io_dat_actv_nz_92,
  input         io_dat_actv_nz_93,
  input         io_dat_actv_nz_94,
  input         io_dat_actv_nz_95,
  input         io_dat_actv_nz_96,
  input         io_dat_actv_nz_97,
  input         io_dat_actv_nz_98,
  input         io_dat_actv_nz_99,
  input         io_dat_actv_nz_100,
  input         io_dat_actv_nz_101,
  input         io_dat_actv_nz_102,
  input         io_dat_actv_nz_103,
  input         io_dat_actv_nz_104,
  input         io_dat_actv_nz_105,
  input         io_dat_actv_nz_106,
  input         io_dat_actv_nz_107,
  input         io_dat_actv_nz_108,
  input         io_dat_actv_nz_109,
  input         io_dat_actv_nz_110,
  input         io_dat_actv_nz_111,
  input         io_dat_actv_nz_112,
  input         io_dat_actv_nz_113,
  input         io_dat_actv_nz_114,
  input         io_dat_actv_nz_115,
  input         io_dat_actv_nz_116,
  input         io_dat_actv_nz_117,
  input         io_dat_actv_nz_118,
  input         io_dat_actv_nz_119,
  input         io_dat_actv_nz_120,
  input         io_dat_actv_nz_121,
  input         io_dat_actv_nz_122,
  input         io_dat_actv_nz_123,
  input         io_dat_actv_nz_124,
  input         io_dat_actv_nz_125,
  input         io_dat_actv_nz_126,
  input         io_dat_actv_nz_127,
  input         io_dat_actv_pvld_0,
  input         io_dat_actv_pvld_1,
  input         io_dat_actv_pvld_2,
  input         io_dat_actv_pvld_3,
  input         io_dat_actv_pvld_4,
  input         io_dat_actv_pvld_5,
  input         io_dat_actv_pvld_6,
  input         io_dat_actv_pvld_7,
  input         io_dat_actv_pvld_8,
  input         io_dat_actv_pvld_9,
  input         io_dat_actv_pvld_10,
  input         io_dat_actv_pvld_11,
  input         io_dat_actv_pvld_12,
  input         io_dat_actv_pvld_13,
  input         io_dat_actv_pvld_14,
  input         io_dat_actv_pvld_15,
  input         io_dat_actv_pvld_16,
  input         io_dat_actv_pvld_17,
  input         io_dat_actv_pvld_18,
  input         io_dat_actv_pvld_19,
  input         io_dat_actv_pvld_20,
  input         io_dat_actv_pvld_21,
  input         io_dat_actv_pvld_22,
  input         io_dat_actv_pvld_23,
  input         io_dat_actv_pvld_24,
  input         io_dat_actv_pvld_25,
  input         io_dat_actv_pvld_26,
  input         io_dat_actv_pvld_27,
  input         io_dat_actv_pvld_28,
  input         io_dat_actv_pvld_29,
  input         io_dat_actv_pvld_30,
  input         io_dat_actv_pvld_31,
  input         io_dat_actv_pvld_32,
  input         io_dat_actv_pvld_33,
  input         io_dat_actv_pvld_34,
  input         io_dat_actv_pvld_35,
  input         io_dat_actv_pvld_36,
  input         io_dat_actv_pvld_37,
  input         io_dat_actv_pvld_38,
  input         io_dat_actv_pvld_39,
  input         io_dat_actv_pvld_40,
  input         io_dat_actv_pvld_41,
  input         io_dat_actv_pvld_42,
  input         io_dat_actv_pvld_43,
  input         io_dat_actv_pvld_44,
  input         io_dat_actv_pvld_45,
  input         io_dat_actv_pvld_46,
  input         io_dat_actv_pvld_47,
  input         io_dat_actv_pvld_48,
  input         io_dat_actv_pvld_49,
  input         io_dat_actv_pvld_50,
  input         io_dat_actv_pvld_51,
  input         io_dat_actv_pvld_52,
  input         io_dat_actv_pvld_53,
  input         io_dat_actv_pvld_54,
  input         io_dat_actv_pvld_55,
  input         io_dat_actv_pvld_56,
  input         io_dat_actv_pvld_57,
  input         io_dat_actv_pvld_58,
  input         io_dat_actv_pvld_59,
  input         io_dat_actv_pvld_60,
  input         io_dat_actv_pvld_61,
  input         io_dat_actv_pvld_62,
  input         io_dat_actv_pvld_63,
  input         io_dat_actv_pvld_64,
  input         io_dat_actv_pvld_65,
  input         io_dat_actv_pvld_66,
  input         io_dat_actv_pvld_67,
  input         io_dat_actv_pvld_68,
  input         io_dat_actv_pvld_69,
  input         io_dat_actv_pvld_70,
  input         io_dat_actv_pvld_71,
  input         io_dat_actv_pvld_72,
  input         io_dat_actv_pvld_73,
  input         io_dat_actv_pvld_74,
  input         io_dat_actv_pvld_75,
  input         io_dat_actv_pvld_76,
  input         io_dat_actv_pvld_77,
  input         io_dat_actv_pvld_78,
  input         io_dat_actv_pvld_79,
  input         io_dat_actv_pvld_80,
  input         io_dat_actv_pvld_81,
  input         io_dat_actv_pvld_82,
  input         io_dat_actv_pvld_83,
  input         io_dat_actv_pvld_84,
  input         io_dat_actv_pvld_85,
  input         io_dat_actv_pvld_86,
  input         io_dat_actv_pvld_87,
  input         io_dat_actv_pvld_88,
  input         io_dat_actv_pvld_89,
  input         io_dat_actv_pvld_90,
  input         io_dat_actv_pvld_91,
  input         io_dat_actv_pvld_92,
  input         io_dat_actv_pvld_93,
  input         io_dat_actv_pvld_94,
  input         io_dat_actv_pvld_95,
  input         io_dat_actv_pvld_96,
  input         io_dat_actv_pvld_97,
  input         io_dat_actv_pvld_98,
  input         io_dat_actv_pvld_99,
  input         io_dat_actv_pvld_100,
  input         io_dat_actv_pvld_101,
  input         io_dat_actv_pvld_102,
  input         io_dat_actv_pvld_103,
  input         io_dat_actv_pvld_104,
  input         io_dat_actv_pvld_105,
  input         io_dat_actv_pvld_106,
  input         io_dat_actv_pvld_107,
  input         io_dat_actv_pvld_108,
  input         io_dat_actv_pvld_109,
  input         io_dat_actv_pvld_110,
  input         io_dat_actv_pvld_111,
  input         io_dat_actv_pvld_112,
  input         io_dat_actv_pvld_113,
  input         io_dat_actv_pvld_114,
  input         io_dat_actv_pvld_115,
  input         io_dat_actv_pvld_116,
  input         io_dat_actv_pvld_117,
  input         io_dat_actv_pvld_118,
  input         io_dat_actv_pvld_119,
  input         io_dat_actv_pvld_120,
  input         io_dat_actv_pvld_121,
  input         io_dat_actv_pvld_122,
  input         io_dat_actv_pvld_123,
  input         io_dat_actv_pvld_124,
  input         io_dat_actv_pvld_125,
  input         io_dat_actv_pvld_126,
  input         io_dat_actv_pvld_127,
  input  [7:0]  io_wt_actv_data_0,
  input  [7:0]  io_wt_actv_data_1,
  input  [7:0]  io_wt_actv_data_2,
  input  [7:0]  io_wt_actv_data_3,
  input  [7:0]  io_wt_actv_data_4,
  input  [7:0]  io_wt_actv_data_5,
  input  [7:0]  io_wt_actv_data_6,
  input  [7:0]  io_wt_actv_data_7,
  input  [7:0]  io_wt_actv_data_8,
  input  [7:0]  io_wt_actv_data_9,
  input  [7:0]  io_wt_actv_data_10,
  input  [7:0]  io_wt_actv_data_11,
  input  [7:0]  io_wt_actv_data_12,
  input  [7:0]  io_wt_actv_data_13,
  input  [7:0]  io_wt_actv_data_14,
  input  [7:0]  io_wt_actv_data_15,
  input  [7:0]  io_wt_actv_data_16,
  input  [7:0]  io_wt_actv_data_17,
  input  [7:0]  io_wt_actv_data_18,
  input  [7:0]  io_wt_actv_data_19,
  input  [7:0]  io_wt_actv_data_20,
  input  [7:0]  io_wt_actv_data_21,
  input  [7:0]  io_wt_actv_data_22,
  input  [7:0]  io_wt_actv_data_23,
  input  [7:0]  io_wt_actv_data_24,
  input  [7:0]  io_wt_actv_data_25,
  input  [7:0]  io_wt_actv_data_26,
  input  [7:0]  io_wt_actv_data_27,
  input  [7:0]  io_wt_actv_data_28,
  input  [7:0]  io_wt_actv_data_29,
  input  [7:0]  io_wt_actv_data_30,
  input  [7:0]  io_wt_actv_data_31,
  input  [7:0]  io_wt_actv_data_32,
  input  [7:0]  io_wt_actv_data_33,
  input  [7:0]  io_wt_actv_data_34,
  input  [7:0]  io_wt_actv_data_35,
  input  [7:0]  io_wt_actv_data_36,
  input  [7:0]  io_wt_actv_data_37,
  input  [7:0]  io_wt_actv_data_38,
  input  [7:0]  io_wt_actv_data_39,
  input  [7:0]  io_wt_actv_data_40,
  input  [7:0]  io_wt_actv_data_41,
  input  [7:0]  io_wt_actv_data_42,
  input  [7:0]  io_wt_actv_data_43,
  input  [7:0]  io_wt_actv_data_44,
  input  [7:0]  io_wt_actv_data_45,
  input  [7:0]  io_wt_actv_data_46,
  input  [7:0]  io_wt_actv_data_47,
  input  [7:0]  io_wt_actv_data_48,
  input  [7:0]  io_wt_actv_data_49,
  input  [7:0]  io_wt_actv_data_50,
  input  [7:0]  io_wt_actv_data_51,
  input  [7:0]  io_wt_actv_data_52,
  input  [7:0]  io_wt_actv_data_53,
  input  [7:0]  io_wt_actv_data_54,
  input  [7:0]  io_wt_actv_data_55,
  input  [7:0]  io_wt_actv_data_56,
  input  [7:0]  io_wt_actv_data_57,
  input  [7:0]  io_wt_actv_data_58,
  input  [7:0]  io_wt_actv_data_59,
  input  [7:0]  io_wt_actv_data_60,
  input  [7:0]  io_wt_actv_data_61,
  input  [7:0]  io_wt_actv_data_62,
  input  [7:0]  io_wt_actv_data_63,
  input  [7:0]  io_wt_actv_data_64,
  input  [7:0]  io_wt_actv_data_65,
  input  [7:0]  io_wt_actv_data_66,
  input  [7:0]  io_wt_actv_data_67,
  input  [7:0]  io_wt_actv_data_68,
  input  [7:0]  io_wt_actv_data_69,
  input  [7:0]  io_wt_actv_data_70,
  input  [7:0]  io_wt_actv_data_71,
  input  [7:0]  io_wt_actv_data_72,
  input  [7:0]  io_wt_actv_data_73,
  input  [7:0]  io_wt_actv_data_74,
  input  [7:0]  io_wt_actv_data_75,
  input  [7:0]  io_wt_actv_data_76,
  input  [7:0]  io_wt_actv_data_77,
  input  [7:0]  io_wt_actv_data_78,
  input  [7:0]  io_wt_actv_data_79,
  input  [7:0]  io_wt_actv_data_80,
  input  [7:0]  io_wt_actv_data_81,
  input  [7:0]  io_wt_actv_data_82,
  input  [7:0]  io_wt_actv_data_83,
  input  [7:0]  io_wt_actv_data_84,
  input  [7:0]  io_wt_actv_data_85,
  input  [7:0]  io_wt_actv_data_86,
  input  [7:0]  io_wt_actv_data_87,
  input  [7:0]  io_wt_actv_data_88,
  input  [7:0]  io_wt_actv_data_89,
  input  [7:0]  io_wt_actv_data_90,
  input  [7:0]  io_wt_actv_data_91,
  input  [7:0]  io_wt_actv_data_92,
  input  [7:0]  io_wt_actv_data_93,
  input  [7:0]  io_wt_actv_data_94,
  input  [7:0]  io_wt_actv_data_95,
  input  [7:0]  io_wt_actv_data_96,
  input  [7:0]  io_wt_actv_data_97,
  input  [7:0]  io_wt_actv_data_98,
  input  [7:0]  io_wt_actv_data_99,
  input  [7:0]  io_wt_actv_data_100,
  input  [7:0]  io_wt_actv_data_101,
  input  [7:0]  io_wt_actv_data_102,
  input  [7:0]  io_wt_actv_data_103,
  input  [7:0]  io_wt_actv_data_104,
  input  [7:0]  io_wt_actv_data_105,
  input  [7:0]  io_wt_actv_data_106,
  input  [7:0]  io_wt_actv_data_107,
  input  [7:0]  io_wt_actv_data_108,
  input  [7:0]  io_wt_actv_data_109,
  input  [7:0]  io_wt_actv_data_110,
  input  [7:0]  io_wt_actv_data_111,
  input  [7:0]  io_wt_actv_data_112,
  input  [7:0]  io_wt_actv_data_113,
  input  [7:0]  io_wt_actv_data_114,
  input  [7:0]  io_wt_actv_data_115,
  input  [7:0]  io_wt_actv_data_116,
  input  [7:0]  io_wt_actv_data_117,
  input  [7:0]  io_wt_actv_data_118,
  input  [7:0]  io_wt_actv_data_119,
  input  [7:0]  io_wt_actv_data_120,
  input  [7:0]  io_wt_actv_data_121,
  input  [7:0]  io_wt_actv_data_122,
  input  [7:0]  io_wt_actv_data_123,
  input  [7:0]  io_wt_actv_data_124,
  input  [7:0]  io_wt_actv_data_125,
  input  [7:0]  io_wt_actv_data_126,
  input  [7:0]  io_wt_actv_data_127,
  input         io_wt_actv_nz_0,
  input         io_wt_actv_nz_1,
  input         io_wt_actv_nz_2,
  input         io_wt_actv_nz_3,
  input         io_wt_actv_nz_4,
  input         io_wt_actv_nz_5,
  input         io_wt_actv_nz_6,
  input         io_wt_actv_nz_7,
  input         io_wt_actv_nz_8,
  input         io_wt_actv_nz_9,
  input         io_wt_actv_nz_10,
  input         io_wt_actv_nz_11,
  input         io_wt_actv_nz_12,
  input         io_wt_actv_nz_13,
  input         io_wt_actv_nz_14,
  input         io_wt_actv_nz_15,
  input         io_wt_actv_nz_16,
  input         io_wt_actv_nz_17,
  input         io_wt_actv_nz_18,
  input         io_wt_actv_nz_19,
  input         io_wt_actv_nz_20,
  input         io_wt_actv_nz_21,
  input         io_wt_actv_nz_22,
  input         io_wt_actv_nz_23,
  input         io_wt_actv_nz_24,
  input         io_wt_actv_nz_25,
  input         io_wt_actv_nz_26,
  input         io_wt_actv_nz_27,
  input         io_wt_actv_nz_28,
  input         io_wt_actv_nz_29,
  input         io_wt_actv_nz_30,
  input         io_wt_actv_nz_31,
  input         io_wt_actv_nz_32,
  input         io_wt_actv_nz_33,
  input         io_wt_actv_nz_34,
  input         io_wt_actv_nz_35,
  input         io_wt_actv_nz_36,
  input         io_wt_actv_nz_37,
  input         io_wt_actv_nz_38,
  input         io_wt_actv_nz_39,
  input         io_wt_actv_nz_40,
  input         io_wt_actv_nz_41,
  input         io_wt_actv_nz_42,
  input         io_wt_actv_nz_43,
  input         io_wt_actv_nz_44,
  input         io_wt_actv_nz_45,
  input         io_wt_actv_nz_46,
  input         io_wt_actv_nz_47,
  input         io_wt_actv_nz_48,
  input         io_wt_actv_nz_49,
  input         io_wt_actv_nz_50,
  input         io_wt_actv_nz_51,
  input         io_wt_actv_nz_52,
  input         io_wt_actv_nz_53,
  input         io_wt_actv_nz_54,
  input         io_wt_actv_nz_55,
  input         io_wt_actv_nz_56,
  input         io_wt_actv_nz_57,
  input         io_wt_actv_nz_58,
  input         io_wt_actv_nz_59,
  input         io_wt_actv_nz_60,
  input         io_wt_actv_nz_61,
  input         io_wt_actv_nz_62,
  input         io_wt_actv_nz_63,
  input         io_wt_actv_nz_64,
  input         io_wt_actv_nz_65,
  input         io_wt_actv_nz_66,
  input         io_wt_actv_nz_67,
  input         io_wt_actv_nz_68,
  input         io_wt_actv_nz_69,
  input         io_wt_actv_nz_70,
  input         io_wt_actv_nz_71,
  input         io_wt_actv_nz_72,
  input         io_wt_actv_nz_73,
  input         io_wt_actv_nz_74,
  input         io_wt_actv_nz_75,
  input         io_wt_actv_nz_76,
  input         io_wt_actv_nz_77,
  input         io_wt_actv_nz_78,
  input         io_wt_actv_nz_79,
  input         io_wt_actv_nz_80,
  input         io_wt_actv_nz_81,
  input         io_wt_actv_nz_82,
  input         io_wt_actv_nz_83,
  input         io_wt_actv_nz_84,
  input         io_wt_actv_nz_85,
  input         io_wt_actv_nz_86,
  input         io_wt_actv_nz_87,
  input         io_wt_actv_nz_88,
  input         io_wt_actv_nz_89,
  input         io_wt_actv_nz_90,
  input         io_wt_actv_nz_91,
  input         io_wt_actv_nz_92,
  input         io_wt_actv_nz_93,
  input         io_wt_actv_nz_94,
  input         io_wt_actv_nz_95,
  input         io_wt_actv_nz_96,
  input         io_wt_actv_nz_97,
  input         io_wt_actv_nz_98,
  input         io_wt_actv_nz_99,
  input         io_wt_actv_nz_100,
  input         io_wt_actv_nz_101,
  input         io_wt_actv_nz_102,
  input         io_wt_actv_nz_103,
  input         io_wt_actv_nz_104,
  input         io_wt_actv_nz_105,
  input         io_wt_actv_nz_106,
  input         io_wt_actv_nz_107,
  input         io_wt_actv_nz_108,
  input         io_wt_actv_nz_109,
  input         io_wt_actv_nz_110,
  input         io_wt_actv_nz_111,
  input         io_wt_actv_nz_112,
  input         io_wt_actv_nz_113,
  input         io_wt_actv_nz_114,
  input         io_wt_actv_nz_115,
  input         io_wt_actv_nz_116,
  input         io_wt_actv_nz_117,
  input         io_wt_actv_nz_118,
  input         io_wt_actv_nz_119,
  input         io_wt_actv_nz_120,
  input         io_wt_actv_nz_121,
  input         io_wt_actv_nz_122,
  input         io_wt_actv_nz_123,
  input         io_wt_actv_nz_124,
  input         io_wt_actv_nz_125,
  input         io_wt_actv_nz_126,
  input         io_wt_actv_nz_127,
  input         io_wt_actv_pvld_0,
  input         io_wt_actv_pvld_1,
  input         io_wt_actv_pvld_2,
  input         io_wt_actv_pvld_3,
  input         io_wt_actv_pvld_4,
  input         io_wt_actv_pvld_5,
  input         io_wt_actv_pvld_6,
  input         io_wt_actv_pvld_7,
  input         io_wt_actv_pvld_8,
  input         io_wt_actv_pvld_9,
  input         io_wt_actv_pvld_10,
  input         io_wt_actv_pvld_11,
  input         io_wt_actv_pvld_12,
  input         io_wt_actv_pvld_13,
  input         io_wt_actv_pvld_14,
  input         io_wt_actv_pvld_15,
  input         io_wt_actv_pvld_16,
  input         io_wt_actv_pvld_17,
  input         io_wt_actv_pvld_18,
  input         io_wt_actv_pvld_19,
  input         io_wt_actv_pvld_20,
  input         io_wt_actv_pvld_21,
  input         io_wt_actv_pvld_22,
  input         io_wt_actv_pvld_23,
  input         io_wt_actv_pvld_24,
  input         io_wt_actv_pvld_25,
  input         io_wt_actv_pvld_26,
  input         io_wt_actv_pvld_27,
  input         io_wt_actv_pvld_28,
  input         io_wt_actv_pvld_29,
  input         io_wt_actv_pvld_30,
  input         io_wt_actv_pvld_31,
  input         io_wt_actv_pvld_32,
  input         io_wt_actv_pvld_33,
  input         io_wt_actv_pvld_34,
  input         io_wt_actv_pvld_35,
  input         io_wt_actv_pvld_36,
  input         io_wt_actv_pvld_37,
  input         io_wt_actv_pvld_38,
  input         io_wt_actv_pvld_39,
  input         io_wt_actv_pvld_40,
  input         io_wt_actv_pvld_41,
  input         io_wt_actv_pvld_42,
  input         io_wt_actv_pvld_43,
  input         io_wt_actv_pvld_44,
  input         io_wt_actv_pvld_45,
  input         io_wt_actv_pvld_46,
  input         io_wt_actv_pvld_47,
  input         io_wt_actv_pvld_48,
  input         io_wt_actv_pvld_49,
  input         io_wt_actv_pvld_50,
  input         io_wt_actv_pvld_51,
  input         io_wt_actv_pvld_52,
  input         io_wt_actv_pvld_53,
  input         io_wt_actv_pvld_54,
  input         io_wt_actv_pvld_55,
  input         io_wt_actv_pvld_56,
  input         io_wt_actv_pvld_57,
  input         io_wt_actv_pvld_58,
  input         io_wt_actv_pvld_59,
  input         io_wt_actv_pvld_60,
  input         io_wt_actv_pvld_61,
  input         io_wt_actv_pvld_62,
  input         io_wt_actv_pvld_63,
  input         io_wt_actv_pvld_64,
  input         io_wt_actv_pvld_65,
  input         io_wt_actv_pvld_66,
  input         io_wt_actv_pvld_67,
  input         io_wt_actv_pvld_68,
  input         io_wt_actv_pvld_69,
  input         io_wt_actv_pvld_70,
  input         io_wt_actv_pvld_71,
  input         io_wt_actv_pvld_72,
  input         io_wt_actv_pvld_73,
  input         io_wt_actv_pvld_74,
  input         io_wt_actv_pvld_75,
  input         io_wt_actv_pvld_76,
  input         io_wt_actv_pvld_77,
  input         io_wt_actv_pvld_78,
  input         io_wt_actv_pvld_79,
  input         io_wt_actv_pvld_80,
  input         io_wt_actv_pvld_81,
  input         io_wt_actv_pvld_82,
  input         io_wt_actv_pvld_83,
  input         io_wt_actv_pvld_84,
  input         io_wt_actv_pvld_85,
  input         io_wt_actv_pvld_86,
  input         io_wt_actv_pvld_87,
  input         io_wt_actv_pvld_88,
  input         io_wt_actv_pvld_89,
  input         io_wt_actv_pvld_90,
  input         io_wt_actv_pvld_91,
  input         io_wt_actv_pvld_92,
  input         io_wt_actv_pvld_93,
  input         io_wt_actv_pvld_94,
  input         io_wt_actv_pvld_95,
  input         io_wt_actv_pvld_96,
  input         io_wt_actv_pvld_97,
  input         io_wt_actv_pvld_98,
  input         io_wt_actv_pvld_99,
  input         io_wt_actv_pvld_100,
  input         io_wt_actv_pvld_101,
  input         io_wt_actv_pvld_102,
  input         io_wt_actv_pvld_103,
  input         io_wt_actv_pvld_104,
  input         io_wt_actv_pvld_105,
  input         io_wt_actv_pvld_106,
  input         io_wt_actv_pvld_107,
  input         io_wt_actv_pvld_108,
  input         io_wt_actv_pvld_109,
  input         io_wt_actv_pvld_110,
  input         io_wt_actv_pvld_111,
  input         io_wt_actv_pvld_112,
  input         io_wt_actv_pvld_113,
  input         io_wt_actv_pvld_114,
  input         io_wt_actv_pvld_115,
  input         io_wt_actv_pvld_116,
  input         io_wt_actv_pvld_117,
  input         io_wt_actv_pvld_118,
  input         io_wt_actv_pvld_119,
  input         io_wt_actv_pvld_120,
  input         io_wt_actv_pvld_121,
  input         io_wt_actv_pvld_122,
  input         io_wt_actv_pvld_123,
  input         io_wt_actv_pvld_124,
  input         io_wt_actv_pvld_125,
  input         io_wt_actv_pvld_126,
  input         io_wt_actv_pvld_127,
  output [22:0] io_mac_out_data,
  output        io_mac_out_pvld
);
  wire  _T_1866; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1867; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1868; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1869; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1871; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1872; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1873; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1874; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_1; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1876; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1877; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1878; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1879; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_2; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1881; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1882; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1883; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1884; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_3; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1886; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1887; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1888; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1889; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_4; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1891; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1892; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1893; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1894; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_5; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1896; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1897; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1898; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1899; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_6; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1901; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1902; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1903; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1904; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_7; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1906; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1907; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1908; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1909; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_8; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1911; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1912; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1913; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1914; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_9; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1916; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1917; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1918; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1919; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_10; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1921; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1922; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1923; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1924; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_11; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1926; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1927; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1928; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1929; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_12; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1931; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1932; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1933; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1934; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_13; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1936; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1937; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1938; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1939; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_14; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1941; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1942; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1943; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1944; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_15; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1946; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1947; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1948; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1949; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_16; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1951; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1952; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1953; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1954; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_17; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1956; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1957; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1958; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1959; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_18; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1961; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1962; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1963; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1964; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_19; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1966; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1967; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1968; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1969; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_20; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1971; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1972; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1973; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1974; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_21; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1976; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1977; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1978; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1979; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_22; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1981; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1982; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1983; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1984; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_23; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1986; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1987; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1988; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1989; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_24; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1991; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1992; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1993; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1994; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_25; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_1996; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_1997; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_1998; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_1999; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_26; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2001; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2002; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2003; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2004; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_27; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2006; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2007; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2008; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2009; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_28; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2011; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2012; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2013; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2014; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_29; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2016; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2017; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2018; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2019; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_30; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2021; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2022; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2023; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2024; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_31; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2026; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2027; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2028; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2029; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_32; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2031; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2032; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2033; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2034; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_33; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2036; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2037; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2038; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2039; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_34; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2041; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2042; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2043; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2044; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_35; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2046; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2047; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2048; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2049; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_36; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2051; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2052; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2053; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2054; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_37; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2056; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2057; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2058; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2059; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_38; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2061; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2062; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2063; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2064; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_39; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2066; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2067; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2068; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2069; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_40; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2071; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2072; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2073; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2074; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_41; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2076; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2077; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2078; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2079; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_42; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2081; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2082; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2083; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2084; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_43; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2086; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2087; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2088; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2089; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_44; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2091; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2092; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2093; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2094; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_45; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2096; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2097; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2098; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2099; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_46; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2101; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2102; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2103; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2104; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_47; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2106; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2107; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2108; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2109; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_48; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2111; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2112; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2113; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2114; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_49; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2116; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2117; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2118; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2119; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_50; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2121; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2122; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2123; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2124; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_51; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2126; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2127; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2128; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2129; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_52; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2131; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2132; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2133; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2134; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_53; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2136; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2137; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2138; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2139; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_54; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2141; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2142; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2143; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2144; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_55; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2146; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2147; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2148; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2149; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_56; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2151; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2152; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2153; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2154; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_57; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2156; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2157; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2158; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2159; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_58; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2161; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2162; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2163; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2164; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_59; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2166; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2167; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2168; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2169; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_60; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2171; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2172; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2173; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2174; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_61; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2176; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2177; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2178; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2179; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_62; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2181; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2182; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2183; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2184; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_63; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2186; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2187; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2188; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2189; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_64; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2191; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2192; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2193; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2194; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_65; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2196; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2197; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2198; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2199; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_66; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2201; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2202; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2203; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2204; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_67; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2206; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2207; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2208; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2209; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_68; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2211; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2212; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2213; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2214; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_69; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2216; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2217; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2218; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2219; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_70; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2221; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2222; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2223; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2224; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_71; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2226; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2227; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2228; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2229; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_72; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2231; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2232; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2233; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2234; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_73; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2236; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2237; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2238; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2239; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_74; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2241; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2242; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2243; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2244; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_75; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2246; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2247; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2248; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2249; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_76; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2251; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2252; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2253; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2254; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_77; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2256; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2257; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2258; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2259; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_78; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2261; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2262; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2263; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2264; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_79; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2266; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2267; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2268; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2269; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_80; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2271; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2272; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2273; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2274; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_81; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2276; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2277; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2278; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2279; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_82; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2281; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2282; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2283; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2284; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_83; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2286; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2287; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2288; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2289; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_84; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2291; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2292; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2293; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2294; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_85; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2296; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2297; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2298; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2299; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_86; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2301; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2302; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2303; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2304; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_87; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2306; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2307; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2308; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2309; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_88; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2311; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2312; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2313; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2314; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_89; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2316; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2317; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2318; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2319; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_90; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2321; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2322; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2323; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2324; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_91; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2326; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2327; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2328; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2329; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_92; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2331; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2332; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2333; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2334; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_93; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2336; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2337; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2338; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2339; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_94; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2341; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2342; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2343; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2344; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_95; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2346; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2347; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2348; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2349; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_96; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2351; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2352; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2353; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2354; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_97; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2356; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2357; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2358; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2359; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_98; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2361; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2362; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2363; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2364; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_99; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2366; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2367; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2368; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2369; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_100; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2371; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2372; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2373; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2374; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_101; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2376; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2377; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2378; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2379; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_102; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2381; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2382; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2383; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2384; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_103; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2386; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2387; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2388; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2389; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_104; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2391; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2392; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2393; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2394; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_105; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2396; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2397; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2398; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2399; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_106; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2401; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2402; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2403; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2404; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_107; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2406; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2407; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2408; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2409; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_108; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2411; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2412; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2413; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2414; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_109; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2416; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2417; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2418; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2419; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_110; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2421; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2422; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2423; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2424; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_111; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2426; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2427; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2428; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2429; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_112; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2431; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2432; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2433; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2434; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_113; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2436; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2437; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2438; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2439; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_114; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2441; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2442; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2443; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2444; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_115; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2446; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2447; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2448; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2449; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_116; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2451; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2452; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2453; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2454; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_117; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2456; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2457; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2458; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2459; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_118; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2461; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2462; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2463; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2464; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_119; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2466; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2467; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2468; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2469; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_120; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2471; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2472; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2473; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2474; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_121; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2476; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2477; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2478; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2479; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_122; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2481; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2482; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2483; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2484; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_123; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2486; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2487; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2488; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2489; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_124; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2491; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2492; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2493; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2494; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_125; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2496; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2497; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2498; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2499; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_126; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire  _T_2501; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  wire  _T_2502; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  wire  _T_2503; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  wire [15:0] _T_2504; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  wire [22:0] _GEN_127; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  wire [15:0] mout_0; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [15:0] mout_1; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [16:0] _T_2506; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_2; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [16:0] _GEN_134; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [17:0] _T_2507; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_3; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [17:0] _GEN_135; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [18:0] _T_2508; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_4; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [18:0] _GEN_136; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [19:0] _T_2509; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_5; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [19:0] _GEN_137; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [20:0] _T_2510; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_6; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [20:0] _GEN_138; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [21:0] _T_2511; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_7; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [21:0] _GEN_139; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [22:0] _T_2512; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_8; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [22:0] _GEN_140; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [23:0] _T_2513; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_9; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [23:0] _GEN_141; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [24:0] _T_2514; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_10; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [24:0] _GEN_142; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [25:0] _T_2515; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_11; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [25:0] _GEN_143; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [26:0] _T_2516; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_12; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [26:0] _GEN_144; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [27:0] _T_2517; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_13; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [27:0] _GEN_145; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [28:0] _T_2518; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_14; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [28:0] _GEN_146; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [29:0] _T_2519; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_15; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [29:0] _GEN_147; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [30:0] _T_2520; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_16; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [30:0] _GEN_148; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [31:0] _T_2521; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_17; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [31:0] _GEN_149; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [32:0] _T_2522; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_18; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [32:0] _GEN_150; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [33:0] _T_2523; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_19; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [33:0] _GEN_151; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [34:0] _T_2524; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_20; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [34:0] _GEN_152; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [35:0] _T_2525; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_21; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [35:0] _GEN_153; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [36:0] _T_2526; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_22; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [36:0] _GEN_154; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [37:0] _T_2527; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_23; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [37:0] _GEN_155; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [38:0] _T_2528; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_24; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [38:0] _GEN_156; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [39:0] _T_2529; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_25; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [39:0] _GEN_157; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [40:0] _T_2530; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_26; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [40:0] _GEN_158; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [41:0] _T_2531; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_27; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [41:0] _GEN_159; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [42:0] _T_2532; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_28; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [42:0] _GEN_160; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [43:0] _T_2533; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_29; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [43:0] _GEN_161; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [44:0] _T_2534; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_30; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [44:0] _GEN_162; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [45:0] _T_2535; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_31; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [45:0] _GEN_163; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [46:0] _T_2536; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_32; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [46:0] _GEN_164; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [47:0] _T_2537; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_33; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [47:0] _GEN_165; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [48:0] _T_2538; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_34; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [48:0] _GEN_166; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [49:0] _T_2539; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_35; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [49:0] _GEN_167; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [50:0] _T_2540; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_36; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [50:0] _GEN_168; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [51:0] _T_2541; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_37; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [51:0] _GEN_169; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [52:0] _T_2542; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_38; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [52:0] _GEN_170; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [53:0] _T_2543; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_39; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [53:0] _GEN_171; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [54:0] _T_2544; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_40; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [54:0] _GEN_172; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [55:0] _T_2545; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_41; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [55:0] _GEN_173; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [56:0] _T_2546; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_42; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [56:0] _GEN_174; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [57:0] _T_2547; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_43; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [57:0] _GEN_175; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [58:0] _T_2548; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_44; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [58:0] _GEN_176; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [59:0] _T_2549; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_45; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [59:0] _GEN_177; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [60:0] _T_2550; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_46; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [60:0] _GEN_178; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [61:0] _T_2551; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_47; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [61:0] _GEN_179; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [62:0] _T_2552; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_48; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [62:0] _GEN_180; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [63:0] _T_2553; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_49; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [63:0] _GEN_181; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [64:0] _T_2554; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_50; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [64:0] _GEN_182; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [65:0] _T_2555; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_51; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [65:0] _GEN_183; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [66:0] _T_2556; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_52; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [66:0] _GEN_184; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [67:0] _T_2557; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_53; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [67:0] _GEN_185; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [68:0] _T_2558; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_54; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [68:0] _GEN_186; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [69:0] _T_2559; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_55; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [69:0] _GEN_187; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [70:0] _T_2560; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_56; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [70:0] _GEN_188; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [71:0] _T_2561; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_57; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [71:0] _GEN_189; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [72:0] _T_2562; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_58; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [72:0] _GEN_190; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [73:0] _T_2563; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_59; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [73:0] _GEN_191; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [74:0] _T_2564; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_60; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [74:0] _GEN_192; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [75:0] _T_2565; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_61; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [75:0] _GEN_193; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [76:0] _T_2566; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_62; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [76:0] _GEN_194; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [77:0] _T_2567; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_63; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [77:0] _GEN_195; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [78:0] _T_2568; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_64; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [78:0] _GEN_196; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [79:0] _T_2569; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_65; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [79:0] _GEN_197; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [80:0] _T_2570; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_66; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [80:0] _GEN_198; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [81:0] _T_2571; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_67; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [81:0] _GEN_199; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [82:0] _T_2572; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_68; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [82:0] _GEN_200; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [83:0] _T_2573; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_69; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [83:0] _GEN_201; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [84:0] _T_2574; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_70; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [84:0] _GEN_202; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [85:0] _T_2575; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_71; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [85:0] _GEN_203; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [86:0] _T_2576; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_72; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [86:0] _GEN_204; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [87:0] _T_2577; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_73; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [87:0] _GEN_205; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [88:0] _T_2578; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_74; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [88:0] _GEN_206; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [89:0] _T_2579; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_75; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [89:0] _GEN_207; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [90:0] _T_2580; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_76; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [90:0] _GEN_208; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [91:0] _T_2581; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_77; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [91:0] _GEN_209; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [92:0] _T_2582; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_78; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [92:0] _GEN_210; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [93:0] _T_2583; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_79; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [93:0] _GEN_211; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [94:0] _T_2584; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_80; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [94:0] _GEN_212; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [95:0] _T_2585; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_81; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [95:0] _GEN_213; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [96:0] _T_2586; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_82; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [96:0] _GEN_214; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [97:0] _T_2587; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_83; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [97:0] _GEN_215; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [98:0] _T_2588; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_84; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [98:0] _GEN_216; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [99:0] _T_2589; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_85; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [99:0] _GEN_217; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [100:0] _T_2590; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_86; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [100:0] _GEN_218; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [101:0] _T_2591; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_87; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [101:0] _GEN_219; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [102:0] _T_2592; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_88; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [102:0] _GEN_220; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [103:0] _T_2593; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_89; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [103:0] _GEN_221; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [104:0] _T_2594; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_90; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [104:0] _GEN_222; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [105:0] _T_2595; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_91; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [105:0] _GEN_223; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [106:0] _T_2596; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_92; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [106:0] _GEN_224; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [107:0] _T_2597; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_93; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [107:0] _GEN_225; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [108:0] _T_2598; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_94; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [108:0] _GEN_226; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [109:0] _T_2599; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_95; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [109:0] _GEN_227; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [110:0] _T_2600; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_96; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [110:0] _GEN_228; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [111:0] _T_2601; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_97; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [111:0] _GEN_229; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [112:0] _T_2602; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_98; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [112:0] _GEN_230; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [113:0] _T_2603; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_99; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [113:0] _GEN_231; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [114:0] _T_2604; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_100; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [114:0] _GEN_232; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [115:0] _T_2605; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_101; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [115:0] _GEN_233; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [116:0] _T_2606; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_102; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [116:0] _GEN_234; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [117:0] _T_2607; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_103; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [117:0] _GEN_235; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [118:0] _T_2608; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_104; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [118:0] _GEN_236; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [119:0] _T_2609; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_105; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [119:0] _GEN_237; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [120:0] _T_2610; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_106; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [120:0] _GEN_238; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [121:0] _T_2611; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_107; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [121:0] _GEN_239; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [122:0] _T_2612; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_108; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [122:0] _GEN_240; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [123:0] _T_2613; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_109; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [123:0] _GEN_241; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [124:0] _T_2614; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_110; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [124:0] _GEN_242; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [125:0] _T_2615; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_111; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [125:0] _GEN_243; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [126:0] _T_2616; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_112; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [126:0] _GEN_244; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [127:0] _T_2617; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_113; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [127:0] _GEN_245; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [128:0] _T_2618; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_114; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [128:0] _GEN_246; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [129:0] _T_2619; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_115; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [129:0] _GEN_247; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [130:0] _T_2620; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_116; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [130:0] _GEN_248; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [131:0] _T_2621; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_117; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [131:0] _GEN_249; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [132:0] _T_2622; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_118; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [132:0] _GEN_250; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [133:0] _T_2623; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_119; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [133:0] _GEN_251; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [134:0] _T_2624; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_120; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [134:0] _GEN_252; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [135:0] _T_2625; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_121; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [135:0] _GEN_253; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [136:0] _T_2626; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_122; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [136:0] _GEN_254; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [137:0] _T_2627; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_123; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [137:0] _GEN_255; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [138:0] _T_2628; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_124; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [138:0] _GEN_256; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [139:0] _T_2629; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_125; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [139:0] _GEN_257; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [140:0] _T_2630; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_126; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [140:0] _GEN_258; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [141:0] _T_2631; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [15:0] mout_127; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  wire [141:0] _GEN_259; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire [142:0] sum_out; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  wire  pp_pvld_d0; // @[NV_NVDLA_CMAC_CORE_mac.scala 62:41]
  reg [142:0] _T_2633; // @[Reg.scala 11:16]
  reg [159:0] _RAND_0;
  reg [142:0] _T_2635; // @[Reg.scala 11:16]
  reg [159:0] _RAND_1;
  reg [142:0] _T_2637; // @[Reg.scala 11:16]
  reg [159:0] _RAND_2;
  reg  _T_2639; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  reg  _T_2641; // @[Reg.scala 11:16]
  reg [31:0] _RAND_4;
  reg  _T_2643; // @[Reg.scala 11:16]
  reg [31:0] _RAND_5;
  assign _T_1866 = io_wt_actv_pvld_0 & io_wt_actv_nz_0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1867 = _T_1866 & io_dat_actv_pvld_0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1868 = _T_1867 & io_dat_actv_nz_0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1869 = io_wt_actv_data_0 * io_dat_actv_data_0; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_0 = _T_1868 ? {{7'd0}, _T_1869} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1871 = io_wt_actv_pvld_1 & io_wt_actv_nz_1; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1872 = _T_1871 & io_dat_actv_pvld_1; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1873 = _T_1872 & io_dat_actv_nz_1; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1874 = io_wt_actv_data_1 * io_dat_actv_data_1; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_1 = _T_1873 ? {{7'd0}, _T_1874} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1876 = io_wt_actv_pvld_2 & io_wt_actv_nz_2; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1877 = _T_1876 & io_dat_actv_pvld_2; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1878 = _T_1877 & io_dat_actv_nz_2; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1879 = io_wt_actv_data_2 * io_dat_actv_data_2; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_2 = _T_1878 ? {{7'd0}, _T_1879} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1881 = io_wt_actv_pvld_3 & io_wt_actv_nz_3; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1882 = _T_1881 & io_dat_actv_pvld_3; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1883 = _T_1882 & io_dat_actv_nz_3; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1884 = io_wt_actv_data_3 * io_dat_actv_data_3; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_3 = _T_1883 ? {{7'd0}, _T_1884} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1886 = io_wt_actv_pvld_4 & io_wt_actv_nz_4; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1887 = _T_1886 & io_dat_actv_pvld_4; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1888 = _T_1887 & io_dat_actv_nz_4; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1889 = io_wt_actv_data_4 * io_dat_actv_data_4; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_4 = _T_1888 ? {{7'd0}, _T_1889} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1891 = io_wt_actv_pvld_5 & io_wt_actv_nz_5; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1892 = _T_1891 & io_dat_actv_pvld_5; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1893 = _T_1892 & io_dat_actv_nz_5; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1894 = io_wt_actv_data_5 * io_dat_actv_data_5; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_5 = _T_1893 ? {{7'd0}, _T_1894} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1896 = io_wt_actv_pvld_6 & io_wt_actv_nz_6; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1897 = _T_1896 & io_dat_actv_pvld_6; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1898 = _T_1897 & io_dat_actv_nz_6; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1899 = io_wt_actv_data_6 * io_dat_actv_data_6; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_6 = _T_1898 ? {{7'd0}, _T_1899} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1901 = io_wt_actv_pvld_7 & io_wt_actv_nz_7; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1902 = _T_1901 & io_dat_actv_pvld_7; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1903 = _T_1902 & io_dat_actv_nz_7; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1904 = io_wt_actv_data_7 * io_dat_actv_data_7; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_7 = _T_1903 ? {{7'd0}, _T_1904} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1906 = io_wt_actv_pvld_8 & io_wt_actv_nz_8; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1907 = _T_1906 & io_dat_actv_pvld_8; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1908 = _T_1907 & io_dat_actv_nz_8; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1909 = io_wt_actv_data_8 * io_dat_actv_data_8; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_8 = _T_1908 ? {{7'd0}, _T_1909} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1911 = io_wt_actv_pvld_9 & io_wt_actv_nz_9; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1912 = _T_1911 & io_dat_actv_pvld_9; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1913 = _T_1912 & io_dat_actv_nz_9; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1914 = io_wt_actv_data_9 * io_dat_actv_data_9; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_9 = _T_1913 ? {{7'd0}, _T_1914} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1916 = io_wt_actv_pvld_10 & io_wt_actv_nz_10; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1917 = _T_1916 & io_dat_actv_pvld_10; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1918 = _T_1917 & io_dat_actv_nz_10; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1919 = io_wt_actv_data_10 * io_dat_actv_data_10; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_10 = _T_1918 ? {{7'd0}, _T_1919} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1921 = io_wt_actv_pvld_11 & io_wt_actv_nz_11; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1922 = _T_1921 & io_dat_actv_pvld_11; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1923 = _T_1922 & io_dat_actv_nz_11; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1924 = io_wt_actv_data_11 * io_dat_actv_data_11; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_11 = _T_1923 ? {{7'd0}, _T_1924} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1926 = io_wt_actv_pvld_12 & io_wt_actv_nz_12; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1927 = _T_1926 & io_dat_actv_pvld_12; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1928 = _T_1927 & io_dat_actv_nz_12; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1929 = io_wt_actv_data_12 * io_dat_actv_data_12; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_12 = _T_1928 ? {{7'd0}, _T_1929} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1931 = io_wt_actv_pvld_13 & io_wt_actv_nz_13; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1932 = _T_1931 & io_dat_actv_pvld_13; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1933 = _T_1932 & io_dat_actv_nz_13; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1934 = io_wt_actv_data_13 * io_dat_actv_data_13; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_13 = _T_1933 ? {{7'd0}, _T_1934} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1936 = io_wt_actv_pvld_14 & io_wt_actv_nz_14; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1937 = _T_1936 & io_dat_actv_pvld_14; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1938 = _T_1937 & io_dat_actv_nz_14; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1939 = io_wt_actv_data_14 * io_dat_actv_data_14; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_14 = _T_1938 ? {{7'd0}, _T_1939} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1941 = io_wt_actv_pvld_15 & io_wt_actv_nz_15; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1942 = _T_1941 & io_dat_actv_pvld_15; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1943 = _T_1942 & io_dat_actv_nz_15; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1944 = io_wt_actv_data_15 * io_dat_actv_data_15; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_15 = _T_1943 ? {{7'd0}, _T_1944} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1946 = io_wt_actv_pvld_16 & io_wt_actv_nz_16; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1947 = _T_1946 & io_dat_actv_pvld_16; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1948 = _T_1947 & io_dat_actv_nz_16; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1949 = io_wt_actv_data_16 * io_dat_actv_data_16; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_16 = _T_1948 ? {{7'd0}, _T_1949} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1951 = io_wt_actv_pvld_17 & io_wt_actv_nz_17; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1952 = _T_1951 & io_dat_actv_pvld_17; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1953 = _T_1952 & io_dat_actv_nz_17; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1954 = io_wt_actv_data_17 * io_dat_actv_data_17; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_17 = _T_1953 ? {{7'd0}, _T_1954} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1956 = io_wt_actv_pvld_18 & io_wt_actv_nz_18; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1957 = _T_1956 & io_dat_actv_pvld_18; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1958 = _T_1957 & io_dat_actv_nz_18; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1959 = io_wt_actv_data_18 * io_dat_actv_data_18; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_18 = _T_1958 ? {{7'd0}, _T_1959} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1961 = io_wt_actv_pvld_19 & io_wt_actv_nz_19; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1962 = _T_1961 & io_dat_actv_pvld_19; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1963 = _T_1962 & io_dat_actv_nz_19; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1964 = io_wt_actv_data_19 * io_dat_actv_data_19; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_19 = _T_1963 ? {{7'd0}, _T_1964} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1966 = io_wt_actv_pvld_20 & io_wt_actv_nz_20; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1967 = _T_1966 & io_dat_actv_pvld_20; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1968 = _T_1967 & io_dat_actv_nz_20; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1969 = io_wt_actv_data_20 * io_dat_actv_data_20; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_20 = _T_1968 ? {{7'd0}, _T_1969} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1971 = io_wt_actv_pvld_21 & io_wt_actv_nz_21; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1972 = _T_1971 & io_dat_actv_pvld_21; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1973 = _T_1972 & io_dat_actv_nz_21; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1974 = io_wt_actv_data_21 * io_dat_actv_data_21; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_21 = _T_1973 ? {{7'd0}, _T_1974} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1976 = io_wt_actv_pvld_22 & io_wt_actv_nz_22; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1977 = _T_1976 & io_dat_actv_pvld_22; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1978 = _T_1977 & io_dat_actv_nz_22; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1979 = io_wt_actv_data_22 * io_dat_actv_data_22; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_22 = _T_1978 ? {{7'd0}, _T_1979} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1981 = io_wt_actv_pvld_23 & io_wt_actv_nz_23; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1982 = _T_1981 & io_dat_actv_pvld_23; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1983 = _T_1982 & io_dat_actv_nz_23; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1984 = io_wt_actv_data_23 * io_dat_actv_data_23; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_23 = _T_1983 ? {{7'd0}, _T_1984} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1986 = io_wt_actv_pvld_24 & io_wt_actv_nz_24; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1987 = _T_1986 & io_dat_actv_pvld_24; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1988 = _T_1987 & io_dat_actv_nz_24; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1989 = io_wt_actv_data_24 * io_dat_actv_data_24; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_24 = _T_1988 ? {{7'd0}, _T_1989} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1991 = io_wt_actv_pvld_25 & io_wt_actv_nz_25; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1992 = _T_1991 & io_dat_actv_pvld_25; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1993 = _T_1992 & io_dat_actv_nz_25; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1994 = io_wt_actv_data_25 * io_dat_actv_data_25; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_25 = _T_1993 ? {{7'd0}, _T_1994} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_1996 = io_wt_actv_pvld_26 & io_wt_actv_nz_26; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_1997 = _T_1996 & io_dat_actv_pvld_26; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_1998 = _T_1997 & io_dat_actv_nz_26; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_1999 = io_wt_actv_data_26 * io_dat_actv_data_26; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_26 = _T_1998 ? {{7'd0}, _T_1999} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2001 = io_wt_actv_pvld_27 & io_wt_actv_nz_27; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2002 = _T_2001 & io_dat_actv_pvld_27; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2003 = _T_2002 & io_dat_actv_nz_27; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2004 = io_wt_actv_data_27 * io_dat_actv_data_27; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_27 = _T_2003 ? {{7'd0}, _T_2004} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2006 = io_wt_actv_pvld_28 & io_wt_actv_nz_28; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2007 = _T_2006 & io_dat_actv_pvld_28; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2008 = _T_2007 & io_dat_actv_nz_28; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2009 = io_wt_actv_data_28 * io_dat_actv_data_28; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_28 = _T_2008 ? {{7'd0}, _T_2009} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2011 = io_wt_actv_pvld_29 & io_wt_actv_nz_29; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2012 = _T_2011 & io_dat_actv_pvld_29; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2013 = _T_2012 & io_dat_actv_nz_29; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2014 = io_wt_actv_data_29 * io_dat_actv_data_29; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_29 = _T_2013 ? {{7'd0}, _T_2014} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2016 = io_wt_actv_pvld_30 & io_wt_actv_nz_30; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2017 = _T_2016 & io_dat_actv_pvld_30; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2018 = _T_2017 & io_dat_actv_nz_30; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2019 = io_wt_actv_data_30 * io_dat_actv_data_30; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_30 = _T_2018 ? {{7'd0}, _T_2019} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2021 = io_wt_actv_pvld_31 & io_wt_actv_nz_31; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2022 = _T_2021 & io_dat_actv_pvld_31; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2023 = _T_2022 & io_dat_actv_nz_31; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2024 = io_wt_actv_data_31 * io_dat_actv_data_31; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_31 = _T_2023 ? {{7'd0}, _T_2024} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2026 = io_wt_actv_pvld_32 & io_wt_actv_nz_32; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2027 = _T_2026 & io_dat_actv_pvld_32; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2028 = _T_2027 & io_dat_actv_nz_32; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2029 = io_wt_actv_data_32 * io_dat_actv_data_32; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_32 = _T_2028 ? {{7'd0}, _T_2029} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2031 = io_wt_actv_pvld_33 & io_wt_actv_nz_33; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2032 = _T_2031 & io_dat_actv_pvld_33; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2033 = _T_2032 & io_dat_actv_nz_33; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2034 = io_wt_actv_data_33 * io_dat_actv_data_33; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_33 = _T_2033 ? {{7'd0}, _T_2034} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2036 = io_wt_actv_pvld_34 & io_wt_actv_nz_34; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2037 = _T_2036 & io_dat_actv_pvld_34; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2038 = _T_2037 & io_dat_actv_nz_34; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2039 = io_wt_actv_data_34 * io_dat_actv_data_34; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_34 = _T_2038 ? {{7'd0}, _T_2039} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2041 = io_wt_actv_pvld_35 & io_wt_actv_nz_35; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2042 = _T_2041 & io_dat_actv_pvld_35; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2043 = _T_2042 & io_dat_actv_nz_35; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2044 = io_wt_actv_data_35 * io_dat_actv_data_35; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_35 = _T_2043 ? {{7'd0}, _T_2044} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2046 = io_wt_actv_pvld_36 & io_wt_actv_nz_36; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2047 = _T_2046 & io_dat_actv_pvld_36; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2048 = _T_2047 & io_dat_actv_nz_36; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2049 = io_wt_actv_data_36 * io_dat_actv_data_36; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_36 = _T_2048 ? {{7'd0}, _T_2049} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2051 = io_wt_actv_pvld_37 & io_wt_actv_nz_37; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2052 = _T_2051 & io_dat_actv_pvld_37; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2053 = _T_2052 & io_dat_actv_nz_37; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2054 = io_wt_actv_data_37 * io_dat_actv_data_37; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_37 = _T_2053 ? {{7'd0}, _T_2054} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2056 = io_wt_actv_pvld_38 & io_wt_actv_nz_38; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2057 = _T_2056 & io_dat_actv_pvld_38; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2058 = _T_2057 & io_dat_actv_nz_38; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2059 = io_wt_actv_data_38 * io_dat_actv_data_38; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_38 = _T_2058 ? {{7'd0}, _T_2059} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2061 = io_wt_actv_pvld_39 & io_wt_actv_nz_39; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2062 = _T_2061 & io_dat_actv_pvld_39; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2063 = _T_2062 & io_dat_actv_nz_39; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2064 = io_wt_actv_data_39 * io_dat_actv_data_39; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_39 = _T_2063 ? {{7'd0}, _T_2064} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2066 = io_wt_actv_pvld_40 & io_wt_actv_nz_40; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2067 = _T_2066 & io_dat_actv_pvld_40; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2068 = _T_2067 & io_dat_actv_nz_40; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2069 = io_wt_actv_data_40 * io_dat_actv_data_40; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_40 = _T_2068 ? {{7'd0}, _T_2069} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2071 = io_wt_actv_pvld_41 & io_wt_actv_nz_41; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2072 = _T_2071 & io_dat_actv_pvld_41; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2073 = _T_2072 & io_dat_actv_nz_41; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2074 = io_wt_actv_data_41 * io_dat_actv_data_41; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_41 = _T_2073 ? {{7'd0}, _T_2074} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2076 = io_wt_actv_pvld_42 & io_wt_actv_nz_42; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2077 = _T_2076 & io_dat_actv_pvld_42; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2078 = _T_2077 & io_dat_actv_nz_42; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2079 = io_wt_actv_data_42 * io_dat_actv_data_42; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_42 = _T_2078 ? {{7'd0}, _T_2079} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2081 = io_wt_actv_pvld_43 & io_wt_actv_nz_43; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2082 = _T_2081 & io_dat_actv_pvld_43; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2083 = _T_2082 & io_dat_actv_nz_43; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2084 = io_wt_actv_data_43 * io_dat_actv_data_43; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_43 = _T_2083 ? {{7'd0}, _T_2084} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2086 = io_wt_actv_pvld_44 & io_wt_actv_nz_44; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2087 = _T_2086 & io_dat_actv_pvld_44; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2088 = _T_2087 & io_dat_actv_nz_44; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2089 = io_wt_actv_data_44 * io_dat_actv_data_44; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_44 = _T_2088 ? {{7'd0}, _T_2089} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2091 = io_wt_actv_pvld_45 & io_wt_actv_nz_45; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2092 = _T_2091 & io_dat_actv_pvld_45; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2093 = _T_2092 & io_dat_actv_nz_45; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2094 = io_wt_actv_data_45 * io_dat_actv_data_45; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_45 = _T_2093 ? {{7'd0}, _T_2094} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2096 = io_wt_actv_pvld_46 & io_wt_actv_nz_46; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2097 = _T_2096 & io_dat_actv_pvld_46; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2098 = _T_2097 & io_dat_actv_nz_46; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2099 = io_wt_actv_data_46 * io_dat_actv_data_46; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_46 = _T_2098 ? {{7'd0}, _T_2099} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2101 = io_wt_actv_pvld_47 & io_wt_actv_nz_47; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2102 = _T_2101 & io_dat_actv_pvld_47; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2103 = _T_2102 & io_dat_actv_nz_47; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2104 = io_wt_actv_data_47 * io_dat_actv_data_47; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_47 = _T_2103 ? {{7'd0}, _T_2104} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2106 = io_wt_actv_pvld_48 & io_wt_actv_nz_48; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2107 = _T_2106 & io_dat_actv_pvld_48; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2108 = _T_2107 & io_dat_actv_nz_48; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2109 = io_wt_actv_data_48 * io_dat_actv_data_48; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_48 = _T_2108 ? {{7'd0}, _T_2109} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2111 = io_wt_actv_pvld_49 & io_wt_actv_nz_49; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2112 = _T_2111 & io_dat_actv_pvld_49; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2113 = _T_2112 & io_dat_actv_nz_49; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2114 = io_wt_actv_data_49 * io_dat_actv_data_49; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_49 = _T_2113 ? {{7'd0}, _T_2114} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2116 = io_wt_actv_pvld_50 & io_wt_actv_nz_50; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2117 = _T_2116 & io_dat_actv_pvld_50; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2118 = _T_2117 & io_dat_actv_nz_50; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2119 = io_wt_actv_data_50 * io_dat_actv_data_50; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_50 = _T_2118 ? {{7'd0}, _T_2119} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2121 = io_wt_actv_pvld_51 & io_wt_actv_nz_51; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2122 = _T_2121 & io_dat_actv_pvld_51; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2123 = _T_2122 & io_dat_actv_nz_51; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2124 = io_wt_actv_data_51 * io_dat_actv_data_51; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_51 = _T_2123 ? {{7'd0}, _T_2124} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2126 = io_wt_actv_pvld_52 & io_wt_actv_nz_52; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2127 = _T_2126 & io_dat_actv_pvld_52; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2128 = _T_2127 & io_dat_actv_nz_52; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2129 = io_wt_actv_data_52 * io_dat_actv_data_52; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_52 = _T_2128 ? {{7'd0}, _T_2129} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2131 = io_wt_actv_pvld_53 & io_wt_actv_nz_53; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2132 = _T_2131 & io_dat_actv_pvld_53; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2133 = _T_2132 & io_dat_actv_nz_53; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2134 = io_wt_actv_data_53 * io_dat_actv_data_53; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_53 = _T_2133 ? {{7'd0}, _T_2134} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2136 = io_wt_actv_pvld_54 & io_wt_actv_nz_54; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2137 = _T_2136 & io_dat_actv_pvld_54; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2138 = _T_2137 & io_dat_actv_nz_54; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2139 = io_wt_actv_data_54 * io_dat_actv_data_54; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_54 = _T_2138 ? {{7'd0}, _T_2139} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2141 = io_wt_actv_pvld_55 & io_wt_actv_nz_55; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2142 = _T_2141 & io_dat_actv_pvld_55; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2143 = _T_2142 & io_dat_actv_nz_55; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2144 = io_wt_actv_data_55 * io_dat_actv_data_55; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_55 = _T_2143 ? {{7'd0}, _T_2144} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2146 = io_wt_actv_pvld_56 & io_wt_actv_nz_56; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2147 = _T_2146 & io_dat_actv_pvld_56; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2148 = _T_2147 & io_dat_actv_nz_56; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2149 = io_wt_actv_data_56 * io_dat_actv_data_56; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_56 = _T_2148 ? {{7'd0}, _T_2149} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2151 = io_wt_actv_pvld_57 & io_wt_actv_nz_57; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2152 = _T_2151 & io_dat_actv_pvld_57; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2153 = _T_2152 & io_dat_actv_nz_57; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2154 = io_wt_actv_data_57 * io_dat_actv_data_57; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_57 = _T_2153 ? {{7'd0}, _T_2154} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2156 = io_wt_actv_pvld_58 & io_wt_actv_nz_58; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2157 = _T_2156 & io_dat_actv_pvld_58; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2158 = _T_2157 & io_dat_actv_nz_58; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2159 = io_wt_actv_data_58 * io_dat_actv_data_58; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_58 = _T_2158 ? {{7'd0}, _T_2159} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2161 = io_wt_actv_pvld_59 & io_wt_actv_nz_59; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2162 = _T_2161 & io_dat_actv_pvld_59; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2163 = _T_2162 & io_dat_actv_nz_59; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2164 = io_wt_actv_data_59 * io_dat_actv_data_59; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_59 = _T_2163 ? {{7'd0}, _T_2164} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2166 = io_wt_actv_pvld_60 & io_wt_actv_nz_60; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2167 = _T_2166 & io_dat_actv_pvld_60; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2168 = _T_2167 & io_dat_actv_nz_60; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2169 = io_wt_actv_data_60 * io_dat_actv_data_60; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_60 = _T_2168 ? {{7'd0}, _T_2169} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2171 = io_wt_actv_pvld_61 & io_wt_actv_nz_61; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2172 = _T_2171 & io_dat_actv_pvld_61; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2173 = _T_2172 & io_dat_actv_nz_61; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2174 = io_wt_actv_data_61 * io_dat_actv_data_61; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_61 = _T_2173 ? {{7'd0}, _T_2174} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2176 = io_wt_actv_pvld_62 & io_wt_actv_nz_62; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2177 = _T_2176 & io_dat_actv_pvld_62; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2178 = _T_2177 & io_dat_actv_nz_62; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2179 = io_wt_actv_data_62 * io_dat_actv_data_62; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_62 = _T_2178 ? {{7'd0}, _T_2179} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2181 = io_wt_actv_pvld_63 & io_wt_actv_nz_63; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2182 = _T_2181 & io_dat_actv_pvld_63; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2183 = _T_2182 & io_dat_actv_nz_63; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2184 = io_wt_actv_data_63 * io_dat_actv_data_63; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_63 = _T_2183 ? {{7'd0}, _T_2184} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2186 = io_wt_actv_pvld_64 & io_wt_actv_nz_64; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2187 = _T_2186 & io_dat_actv_pvld_64; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2188 = _T_2187 & io_dat_actv_nz_64; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2189 = io_wt_actv_data_64 * io_dat_actv_data_64; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_64 = _T_2188 ? {{7'd0}, _T_2189} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2191 = io_wt_actv_pvld_65 & io_wt_actv_nz_65; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2192 = _T_2191 & io_dat_actv_pvld_65; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2193 = _T_2192 & io_dat_actv_nz_65; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2194 = io_wt_actv_data_65 * io_dat_actv_data_65; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_65 = _T_2193 ? {{7'd0}, _T_2194} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2196 = io_wt_actv_pvld_66 & io_wt_actv_nz_66; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2197 = _T_2196 & io_dat_actv_pvld_66; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2198 = _T_2197 & io_dat_actv_nz_66; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2199 = io_wt_actv_data_66 * io_dat_actv_data_66; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_66 = _T_2198 ? {{7'd0}, _T_2199} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2201 = io_wt_actv_pvld_67 & io_wt_actv_nz_67; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2202 = _T_2201 & io_dat_actv_pvld_67; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2203 = _T_2202 & io_dat_actv_nz_67; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2204 = io_wt_actv_data_67 * io_dat_actv_data_67; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_67 = _T_2203 ? {{7'd0}, _T_2204} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2206 = io_wt_actv_pvld_68 & io_wt_actv_nz_68; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2207 = _T_2206 & io_dat_actv_pvld_68; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2208 = _T_2207 & io_dat_actv_nz_68; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2209 = io_wt_actv_data_68 * io_dat_actv_data_68; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_68 = _T_2208 ? {{7'd0}, _T_2209} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2211 = io_wt_actv_pvld_69 & io_wt_actv_nz_69; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2212 = _T_2211 & io_dat_actv_pvld_69; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2213 = _T_2212 & io_dat_actv_nz_69; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2214 = io_wt_actv_data_69 * io_dat_actv_data_69; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_69 = _T_2213 ? {{7'd0}, _T_2214} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2216 = io_wt_actv_pvld_70 & io_wt_actv_nz_70; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2217 = _T_2216 & io_dat_actv_pvld_70; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2218 = _T_2217 & io_dat_actv_nz_70; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2219 = io_wt_actv_data_70 * io_dat_actv_data_70; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_70 = _T_2218 ? {{7'd0}, _T_2219} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2221 = io_wt_actv_pvld_71 & io_wt_actv_nz_71; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2222 = _T_2221 & io_dat_actv_pvld_71; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2223 = _T_2222 & io_dat_actv_nz_71; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2224 = io_wt_actv_data_71 * io_dat_actv_data_71; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_71 = _T_2223 ? {{7'd0}, _T_2224} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2226 = io_wt_actv_pvld_72 & io_wt_actv_nz_72; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2227 = _T_2226 & io_dat_actv_pvld_72; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2228 = _T_2227 & io_dat_actv_nz_72; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2229 = io_wt_actv_data_72 * io_dat_actv_data_72; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_72 = _T_2228 ? {{7'd0}, _T_2229} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2231 = io_wt_actv_pvld_73 & io_wt_actv_nz_73; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2232 = _T_2231 & io_dat_actv_pvld_73; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2233 = _T_2232 & io_dat_actv_nz_73; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2234 = io_wt_actv_data_73 * io_dat_actv_data_73; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_73 = _T_2233 ? {{7'd0}, _T_2234} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2236 = io_wt_actv_pvld_74 & io_wt_actv_nz_74; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2237 = _T_2236 & io_dat_actv_pvld_74; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2238 = _T_2237 & io_dat_actv_nz_74; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2239 = io_wt_actv_data_74 * io_dat_actv_data_74; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_74 = _T_2238 ? {{7'd0}, _T_2239} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2241 = io_wt_actv_pvld_75 & io_wt_actv_nz_75; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2242 = _T_2241 & io_dat_actv_pvld_75; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2243 = _T_2242 & io_dat_actv_nz_75; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2244 = io_wt_actv_data_75 * io_dat_actv_data_75; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_75 = _T_2243 ? {{7'd0}, _T_2244} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2246 = io_wt_actv_pvld_76 & io_wt_actv_nz_76; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2247 = _T_2246 & io_dat_actv_pvld_76; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2248 = _T_2247 & io_dat_actv_nz_76; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2249 = io_wt_actv_data_76 * io_dat_actv_data_76; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_76 = _T_2248 ? {{7'd0}, _T_2249} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2251 = io_wt_actv_pvld_77 & io_wt_actv_nz_77; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2252 = _T_2251 & io_dat_actv_pvld_77; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2253 = _T_2252 & io_dat_actv_nz_77; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2254 = io_wt_actv_data_77 * io_dat_actv_data_77; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_77 = _T_2253 ? {{7'd0}, _T_2254} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2256 = io_wt_actv_pvld_78 & io_wt_actv_nz_78; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2257 = _T_2256 & io_dat_actv_pvld_78; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2258 = _T_2257 & io_dat_actv_nz_78; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2259 = io_wt_actv_data_78 * io_dat_actv_data_78; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_78 = _T_2258 ? {{7'd0}, _T_2259} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2261 = io_wt_actv_pvld_79 & io_wt_actv_nz_79; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2262 = _T_2261 & io_dat_actv_pvld_79; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2263 = _T_2262 & io_dat_actv_nz_79; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2264 = io_wt_actv_data_79 * io_dat_actv_data_79; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_79 = _T_2263 ? {{7'd0}, _T_2264} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2266 = io_wt_actv_pvld_80 & io_wt_actv_nz_80; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2267 = _T_2266 & io_dat_actv_pvld_80; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2268 = _T_2267 & io_dat_actv_nz_80; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2269 = io_wt_actv_data_80 * io_dat_actv_data_80; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_80 = _T_2268 ? {{7'd0}, _T_2269} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2271 = io_wt_actv_pvld_81 & io_wt_actv_nz_81; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2272 = _T_2271 & io_dat_actv_pvld_81; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2273 = _T_2272 & io_dat_actv_nz_81; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2274 = io_wt_actv_data_81 * io_dat_actv_data_81; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_81 = _T_2273 ? {{7'd0}, _T_2274} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2276 = io_wt_actv_pvld_82 & io_wt_actv_nz_82; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2277 = _T_2276 & io_dat_actv_pvld_82; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2278 = _T_2277 & io_dat_actv_nz_82; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2279 = io_wt_actv_data_82 * io_dat_actv_data_82; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_82 = _T_2278 ? {{7'd0}, _T_2279} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2281 = io_wt_actv_pvld_83 & io_wt_actv_nz_83; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2282 = _T_2281 & io_dat_actv_pvld_83; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2283 = _T_2282 & io_dat_actv_nz_83; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2284 = io_wt_actv_data_83 * io_dat_actv_data_83; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_83 = _T_2283 ? {{7'd0}, _T_2284} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2286 = io_wt_actv_pvld_84 & io_wt_actv_nz_84; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2287 = _T_2286 & io_dat_actv_pvld_84; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2288 = _T_2287 & io_dat_actv_nz_84; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2289 = io_wt_actv_data_84 * io_dat_actv_data_84; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_84 = _T_2288 ? {{7'd0}, _T_2289} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2291 = io_wt_actv_pvld_85 & io_wt_actv_nz_85; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2292 = _T_2291 & io_dat_actv_pvld_85; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2293 = _T_2292 & io_dat_actv_nz_85; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2294 = io_wt_actv_data_85 * io_dat_actv_data_85; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_85 = _T_2293 ? {{7'd0}, _T_2294} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2296 = io_wt_actv_pvld_86 & io_wt_actv_nz_86; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2297 = _T_2296 & io_dat_actv_pvld_86; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2298 = _T_2297 & io_dat_actv_nz_86; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2299 = io_wt_actv_data_86 * io_dat_actv_data_86; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_86 = _T_2298 ? {{7'd0}, _T_2299} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2301 = io_wt_actv_pvld_87 & io_wt_actv_nz_87; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2302 = _T_2301 & io_dat_actv_pvld_87; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2303 = _T_2302 & io_dat_actv_nz_87; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2304 = io_wt_actv_data_87 * io_dat_actv_data_87; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_87 = _T_2303 ? {{7'd0}, _T_2304} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2306 = io_wt_actv_pvld_88 & io_wt_actv_nz_88; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2307 = _T_2306 & io_dat_actv_pvld_88; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2308 = _T_2307 & io_dat_actv_nz_88; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2309 = io_wt_actv_data_88 * io_dat_actv_data_88; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_88 = _T_2308 ? {{7'd0}, _T_2309} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2311 = io_wt_actv_pvld_89 & io_wt_actv_nz_89; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2312 = _T_2311 & io_dat_actv_pvld_89; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2313 = _T_2312 & io_dat_actv_nz_89; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2314 = io_wt_actv_data_89 * io_dat_actv_data_89; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_89 = _T_2313 ? {{7'd0}, _T_2314} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2316 = io_wt_actv_pvld_90 & io_wt_actv_nz_90; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2317 = _T_2316 & io_dat_actv_pvld_90; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2318 = _T_2317 & io_dat_actv_nz_90; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2319 = io_wt_actv_data_90 * io_dat_actv_data_90; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_90 = _T_2318 ? {{7'd0}, _T_2319} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2321 = io_wt_actv_pvld_91 & io_wt_actv_nz_91; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2322 = _T_2321 & io_dat_actv_pvld_91; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2323 = _T_2322 & io_dat_actv_nz_91; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2324 = io_wt_actv_data_91 * io_dat_actv_data_91; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_91 = _T_2323 ? {{7'd0}, _T_2324} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2326 = io_wt_actv_pvld_92 & io_wt_actv_nz_92; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2327 = _T_2326 & io_dat_actv_pvld_92; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2328 = _T_2327 & io_dat_actv_nz_92; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2329 = io_wt_actv_data_92 * io_dat_actv_data_92; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_92 = _T_2328 ? {{7'd0}, _T_2329} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2331 = io_wt_actv_pvld_93 & io_wt_actv_nz_93; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2332 = _T_2331 & io_dat_actv_pvld_93; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2333 = _T_2332 & io_dat_actv_nz_93; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2334 = io_wt_actv_data_93 * io_dat_actv_data_93; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_93 = _T_2333 ? {{7'd0}, _T_2334} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2336 = io_wt_actv_pvld_94 & io_wt_actv_nz_94; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2337 = _T_2336 & io_dat_actv_pvld_94; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2338 = _T_2337 & io_dat_actv_nz_94; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2339 = io_wt_actv_data_94 * io_dat_actv_data_94; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_94 = _T_2338 ? {{7'd0}, _T_2339} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2341 = io_wt_actv_pvld_95 & io_wt_actv_nz_95; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2342 = _T_2341 & io_dat_actv_pvld_95; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2343 = _T_2342 & io_dat_actv_nz_95; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2344 = io_wt_actv_data_95 * io_dat_actv_data_95; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_95 = _T_2343 ? {{7'd0}, _T_2344} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2346 = io_wt_actv_pvld_96 & io_wt_actv_nz_96; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2347 = _T_2346 & io_dat_actv_pvld_96; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2348 = _T_2347 & io_dat_actv_nz_96; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2349 = io_wt_actv_data_96 * io_dat_actv_data_96; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_96 = _T_2348 ? {{7'd0}, _T_2349} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2351 = io_wt_actv_pvld_97 & io_wt_actv_nz_97; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2352 = _T_2351 & io_dat_actv_pvld_97; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2353 = _T_2352 & io_dat_actv_nz_97; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2354 = io_wt_actv_data_97 * io_dat_actv_data_97; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_97 = _T_2353 ? {{7'd0}, _T_2354} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2356 = io_wt_actv_pvld_98 & io_wt_actv_nz_98; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2357 = _T_2356 & io_dat_actv_pvld_98; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2358 = _T_2357 & io_dat_actv_nz_98; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2359 = io_wt_actv_data_98 * io_dat_actv_data_98; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_98 = _T_2358 ? {{7'd0}, _T_2359} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2361 = io_wt_actv_pvld_99 & io_wt_actv_nz_99; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2362 = _T_2361 & io_dat_actv_pvld_99; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2363 = _T_2362 & io_dat_actv_nz_99; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2364 = io_wt_actv_data_99 * io_dat_actv_data_99; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_99 = _T_2363 ? {{7'd0}, _T_2364} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2366 = io_wt_actv_pvld_100 & io_wt_actv_nz_100; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2367 = _T_2366 & io_dat_actv_pvld_100; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2368 = _T_2367 & io_dat_actv_nz_100; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2369 = io_wt_actv_data_100 * io_dat_actv_data_100; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_100 = _T_2368 ? {{7'd0}, _T_2369} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2371 = io_wt_actv_pvld_101 & io_wt_actv_nz_101; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2372 = _T_2371 & io_dat_actv_pvld_101; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2373 = _T_2372 & io_dat_actv_nz_101; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2374 = io_wt_actv_data_101 * io_dat_actv_data_101; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_101 = _T_2373 ? {{7'd0}, _T_2374} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2376 = io_wt_actv_pvld_102 & io_wt_actv_nz_102; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2377 = _T_2376 & io_dat_actv_pvld_102; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2378 = _T_2377 & io_dat_actv_nz_102; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2379 = io_wt_actv_data_102 * io_dat_actv_data_102; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_102 = _T_2378 ? {{7'd0}, _T_2379} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2381 = io_wt_actv_pvld_103 & io_wt_actv_nz_103; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2382 = _T_2381 & io_dat_actv_pvld_103; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2383 = _T_2382 & io_dat_actv_nz_103; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2384 = io_wt_actv_data_103 * io_dat_actv_data_103; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_103 = _T_2383 ? {{7'd0}, _T_2384} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2386 = io_wt_actv_pvld_104 & io_wt_actv_nz_104; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2387 = _T_2386 & io_dat_actv_pvld_104; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2388 = _T_2387 & io_dat_actv_nz_104; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2389 = io_wt_actv_data_104 * io_dat_actv_data_104; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_104 = _T_2388 ? {{7'd0}, _T_2389} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2391 = io_wt_actv_pvld_105 & io_wt_actv_nz_105; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2392 = _T_2391 & io_dat_actv_pvld_105; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2393 = _T_2392 & io_dat_actv_nz_105; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2394 = io_wt_actv_data_105 * io_dat_actv_data_105; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_105 = _T_2393 ? {{7'd0}, _T_2394} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2396 = io_wt_actv_pvld_106 & io_wt_actv_nz_106; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2397 = _T_2396 & io_dat_actv_pvld_106; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2398 = _T_2397 & io_dat_actv_nz_106; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2399 = io_wt_actv_data_106 * io_dat_actv_data_106; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_106 = _T_2398 ? {{7'd0}, _T_2399} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2401 = io_wt_actv_pvld_107 & io_wt_actv_nz_107; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2402 = _T_2401 & io_dat_actv_pvld_107; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2403 = _T_2402 & io_dat_actv_nz_107; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2404 = io_wt_actv_data_107 * io_dat_actv_data_107; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_107 = _T_2403 ? {{7'd0}, _T_2404} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2406 = io_wt_actv_pvld_108 & io_wt_actv_nz_108; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2407 = _T_2406 & io_dat_actv_pvld_108; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2408 = _T_2407 & io_dat_actv_nz_108; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2409 = io_wt_actv_data_108 * io_dat_actv_data_108; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_108 = _T_2408 ? {{7'd0}, _T_2409} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2411 = io_wt_actv_pvld_109 & io_wt_actv_nz_109; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2412 = _T_2411 & io_dat_actv_pvld_109; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2413 = _T_2412 & io_dat_actv_nz_109; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2414 = io_wt_actv_data_109 * io_dat_actv_data_109; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_109 = _T_2413 ? {{7'd0}, _T_2414} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2416 = io_wt_actv_pvld_110 & io_wt_actv_nz_110; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2417 = _T_2416 & io_dat_actv_pvld_110; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2418 = _T_2417 & io_dat_actv_nz_110; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2419 = io_wt_actv_data_110 * io_dat_actv_data_110; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_110 = _T_2418 ? {{7'd0}, _T_2419} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2421 = io_wt_actv_pvld_111 & io_wt_actv_nz_111; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2422 = _T_2421 & io_dat_actv_pvld_111; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2423 = _T_2422 & io_dat_actv_nz_111; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2424 = io_wt_actv_data_111 * io_dat_actv_data_111; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_111 = _T_2423 ? {{7'd0}, _T_2424} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2426 = io_wt_actv_pvld_112 & io_wt_actv_nz_112; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2427 = _T_2426 & io_dat_actv_pvld_112; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2428 = _T_2427 & io_dat_actv_nz_112; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2429 = io_wt_actv_data_112 * io_dat_actv_data_112; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_112 = _T_2428 ? {{7'd0}, _T_2429} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2431 = io_wt_actv_pvld_113 & io_wt_actv_nz_113; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2432 = _T_2431 & io_dat_actv_pvld_113; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2433 = _T_2432 & io_dat_actv_nz_113; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2434 = io_wt_actv_data_113 * io_dat_actv_data_113; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_113 = _T_2433 ? {{7'd0}, _T_2434} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2436 = io_wt_actv_pvld_114 & io_wt_actv_nz_114; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2437 = _T_2436 & io_dat_actv_pvld_114; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2438 = _T_2437 & io_dat_actv_nz_114; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2439 = io_wt_actv_data_114 * io_dat_actv_data_114; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_114 = _T_2438 ? {{7'd0}, _T_2439} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2441 = io_wt_actv_pvld_115 & io_wt_actv_nz_115; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2442 = _T_2441 & io_dat_actv_pvld_115; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2443 = _T_2442 & io_dat_actv_nz_115; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2444 = io_wt_actv_data_115 * io_dat_actv_data_115; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_115 = _T_2443 ? {{7'd0}, _T_2444} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2446 = io_wt_actv_pvld_116 & io_wt_actv_nz_116; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2447 = _T_2446 & io_dat_actv_pvld_116; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2448 = _T_2447 & io_dat_actv_nz_116; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2449 = io_wt_actv_data_116 * io_dat_actv_data_116; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_116 = _T_2448 ? {{7'd0}, _T_2449} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2451 = io_wt_actv_pvld_117 & io_wt_actv_nz_117; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2452 = _T_2451 & io_dat_actv_pvld_117; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2453 = _T_2452 & io_dat_actv_nz_117; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2454 = io_wt_actv_data_117 * io_dat_actv_data_117; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_117 = _T_2453 ? {{7'd0}, _T_2454} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2456 = io_wt_actv_pvld_118 & io_wt_actv_nz_118; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2457 = _T_2456 & io_dat_actv_pvld_118; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2458 = _T_2457 & io_dat_actv_nz_118; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2459 = io_wt_actv_data_118 * io_dat_actv_data_118; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_118 = _T_2458 ? {{7'd0}, _T_2459} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2461 = io_wt_actv_pvld_119 & io_wt_actv_nz_119; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2462 = _T_2461 & io_dat_actv_pvld_119; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2463 = _T_2462 & io_dat_actv_nz_119; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2464 = io_wt_actv_data_119 * io_dat_actv_data_119; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_119 = _T_2463 ? {{7'd0}, _T_2464} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2466 = io_wt_actv_pvld_120 & io_wt_actv_nz_120; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2467 = _T_2466 & io_dat_actv_pvld_120; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2468 = _T_2467 & io_dat_actv_nz_120; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2469 = io_wt_actv_data_120 * io_dat_actv_data_120; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_120 = _T_2468 ? {{7'd0}, _T_2469} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2471 = io_wt_actv_pvld_121 & io_wt_actv_nz_121; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2472 = _T_2471 & io_dat_actv_pvld_121; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2473 = _T_2472 & io_dat_actv_nz_121; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2474 = io_wt_actv_data_121 * io_dat_actv_data_121; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_121 = _T_2473 ? {{7'd0}, _T_2474} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2476 = io_wt_actv_pvld_122 & io_wt_actv_nz_122; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2477 = _T_2476 & io_dat_actv_pvld_122; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2478 = _T_2477 & io_dat_actv_nz_122; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2479 = io_wt_actv_data_122 * io_dat_actv_data_122; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_122 = _T_2478 ? {{7'd0}, _T_2479} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2481 = io_wt_actv_pvld_123 & io_wt_actv_nz_123; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2482 = _T_2481 & io_dat_actv_pvld_123; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2483 = _T_2482 & io_dat_actv_nz_123; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2484 = io_wt_actv_data_123 * io_dat_actv_data_123; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_123 = _T_2483 ? {{7'd0}, _T_2484} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2486 = io_wt_actv_pvld_124 & io_wt_actv_nz_124; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2487 = _T_2486 & io_dat_actv_pvld_124; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2488 = _T_2487 & io_dat_actv_nz_124; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2489 = io_wt_actv_data_124 * io_dat_actv_data_124; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_124 = _T_2488 ? {{7'd0}, _T_2489} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2491 = io_wt_actv_pvld_125 & io_wt_actv_nz_125; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2492 = _T_2491 & io_dat_actv_pvld_125; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2493 = _T_2492 & io_dat_actv_nz_125; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2494 = io_wt_actv_data_125 * io_dat_actv_data_125; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_125 = _T_2493 ? {{7'd0}, _T_2494} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2496 = io_wt_actv_pvld_126 & io_wt_actv_nz_126; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2497 = _T_2496 & io_dat_actv_pvld_126; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2498 = _T_2497 & io_dat_actv_nz_126; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2499 = io_wt_actv_data_126 * io_dat_actv_data_126; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_126 = _T_2498 ? {{7'd0}, _T_2499} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign _T_2501 = io_wt_actv_pvld_127 & io_wt_actv_nz_127; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:32]
  assign _T_2502 = _T_2501 & io_dat_actv_pvld_127; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:49]
  assign _T_2503 = _T_2502 & io_dat_actv_nz_127; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:69]
  assign _T_2504 = io_wt_actv_data_127 * io_dat_actv_data_127; // @[NV_NVDLA_CMAC_CORE_mac.scala 52:43]
  assign _GEN_127 = _T_2503 ? {{7'd0}, _T_2504} : 23'h0; // @[NV_NVDLA_CMAC_CORE_mac.scala 51:88]
  assign mout_0 = _GEN_0[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign mout_1 = _GEN_1[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _T_2506 = mout_0 + mout_1; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_2 = _GEN_2[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_134 = {{1'd0}, mout_2}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2507 = _T_2506 + _GEN_134; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_3 = _GEN_3[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_135 = {{2'd0}, mout_3}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2508 = _T_2507 + _GEN_135; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_4 = _GEN_4[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_136 = {{3'd0}, mout_4}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2509 = _T_2508 + _GEN_136; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_5 = _GEN_5[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_137 = {{4'd0}, mout_5}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2510 = _T_2509 + _GEN_137; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_6 = _GEN_6[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_138 = {{5'd0}, mout_6}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2511 = _T_2510 + _GEN_138; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_7 = _GEN_7[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_139 = {{6'd0}, mout_7}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2512 = _T_2511 + _GEN_139; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_8 = _GEN_8[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_140 = {{7'd0}, mout_8}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2513 = _T_2512 + _GEN_140; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_9 = _GEN_9[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_141 = {{8'd0}, mout_9}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2514 = _T_2513 + _GEN_141; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_10 = _GEN_10[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_142 = {{9'd0}, mout_10}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2515 = _T_2514 + _GEN_142; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_11 = _GEN_11[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_143 = {{10'd0}, mout_11}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2516 = _T_2515 + _GEN_143; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_12 = _GEN_12[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_144 = {{11'd0}, mout_12}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2517 = _T_2516 + _GEN_144; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_13 = _GEN_13[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_145 = {{12'd0}, mout_13}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2518 = _T_2517 + _GEN_145; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_14 = _GEN_14[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_146 = {{13'd0}, mout_14}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2519 = _T_2518 + _GEN_146; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_15 = _GEN_15[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_147 = {{14'd0}, mout_15}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2520 = _T_2519 + _GEN_147; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_16 = _GEN_16[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_148 = {{15'd0}, mout_16}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2521 = _T_2520 + _GEN_148; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_17 = _GEN_17[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_149 = {{16'd0}, mout_17}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2522 = _T_2521 + _GEN_149; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_18 = _GEN_18[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_150 = {{17'd0}, mout_18}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2523 = _T_2522 + _GEN_150; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_19 = _GEN_19[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_151 = {{18'd0}, mout_19}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2524 = _T_2523 + _GEN_151; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_20 = _GEN_20[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_152 = {{19'd0}, mout_20}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2525 = _T_2524 + _GEN_152; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_21 = _GEN_21[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_153 = {{20'd0}, mout_21}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2526 = _T_2525 + _GEN_153; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_22 = _GEN_22[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_154 = {{21'd0}, mout_22}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2527 = _T_2526 + _GEN_154; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_23 = _GEN_23[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_155 = {{22'd0}, mout_23}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2528 = _T_2527 + _GEN_155; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_24 = _GEN_24[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_156 = {{23'd0}, mout_24}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2529 = _T_2528 + _GEN_156; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_25 = _GEN_25[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_157 = {{24'd0}, mout_25}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2530 = _T_2529 + _GEN_157; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_26 = _GEN_26[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_158 = {{25'd0}, mout_26}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2531 = _T_2530 + _GEN_158; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_27 = _GEN_27[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_159 = {{26'd0}, mout_27}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2532 = _T_2531 + _GEN_159; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_28 = _GEN_28[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_160 = {{27'd0}, mout_28}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2533 = _T_2532 + _GEN_160; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_29 = _GEN_29[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_161 = {{28'd0}, mout_29}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2534 = _T_2533 + _GEN_161; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_30 = _GEN_30[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_162 = {{29'd0}, mout_30}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2535 = _T_2534 + _GEN_162; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_31 = _GEN_31[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_163 = {{30'd0}, mout_31}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2536 = _T_2535 + _GEN_163; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_32 = _GEN_32[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_164 = {{31'd0}, mout_32}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2537 = _T_2536 + _GEN_164; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_33 = _GEN_33[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_165 = {{32'd0}, mout_33}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2538 = _T_2537 + _GEN_165; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_34 = _GEN_34[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_166 = {{33'd0}, mout_34}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2539 = _T_2538 + _GEN_166; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_35 = _GEN_35[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_167 = {{34'd0}, mout_35}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2540 = _T_2539 + _GEN_167; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_36 = _GEN_36[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_168 = {{35'd0}, mout_36}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2541 = _T_2540 + _GEN_168; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_37 = _GEN_37[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_169 = {{36'd0}, mout_37}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2542 = _T_2541 + _GEN_169; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_38 = _GEN_38[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_170 = {{37'd0}, mout_38}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2543 = _T_2542 + _GEN_170; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_39 = _GEN_39[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_171 = {{38'd0}, mout_39}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2544 = _T_2543 + _GEN_171; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_40 = _GEN_40[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_172 = {{39'd0}, mout_40}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2545 = _T_2544 + _GEN_172; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_41 = _GEN_41[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_173 = {{40'd0}, mout_41}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2546 = _T_2545 + _GEN_173; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_42 = _GEN_42[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_174 = {{41'd0}, mout_42}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2547 = _T_2546 + _GEN_174; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_43 = _GEN_43[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_175 = {{42'd0}, mout_43}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2548 = _T_2547 + _GEN_175; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_44 = _GEN_44[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_176 = {{43'd0}, mout_44}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2549 = _T_2548 + _GEN_176; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_45 = _GEN_45[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_177 = {{44'd0}, mout_45}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2550 = _T_2549 + _GEN_177; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_46 = _GEN_46[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_178 = {{45'd0}, mout_46}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2551 = _T_2550 + _GEN_178; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_47 = _GEN_47[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_179 = {{46'd0}, mout_47}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2552 = _T_2551 + _GEN_179; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_48 = _GEN_48[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_180 = {{47'd0}, mout_48}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2553 = _T_2552 + _GEN_180; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_49 = _GEN_49[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_181 = {{48'd0}, mout_49}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2554 = _T_2553 + _GEN_181; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_50 = _GEN_50[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_182 = {{49'd0}, mout_50}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2555 = _T_2554 + _GEN_182; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_51 = _GEN_51[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_183 = {{50'd0}, mout_51}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2556 = _T_2555 + _GEN_183; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_52 = _GEN_52[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_184 = {{51'd0}, mout_52}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2557 = _T_2556 + _GEN_184; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_53 = _GEN_53[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_185 = {{52'd0}, mout_53}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2558 = _T_2557 + _GEN_185; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_54 = _GEN_54[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_186 = {{53'd0}, mout_54}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2559 = _T_2558 + _GEN_186; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_55 = _GEN_55[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_187 = {{54'd0}, mout_55}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2560 = _T_2559 + _GEN_187; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_56 = _GEN_56[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_188 = {{55'd0}, mout_56}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2561 = _T_2560 + _GEN_188; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_57 = _GEN_57[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_189 = {{56'd0}, mout_57}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2562 = _T_2561 + _GEN_189; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_58 = _GEN_58[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_190 = {{57'd0}, mout_58}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2563 = _T_2562 + _GEN_190; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_59 = _GEN_59[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_191 = {{58'd0}, mout_59}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2564 = _T_2563 + _GEN_191; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_60 = _GEN_60[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_192 = {{59'd0}, mout_60}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2565 = _T_2564 + _GEN_192; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_61 = _GEN_61[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_193 = {{60'd0}, mout_61}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2566 = _T_2565 + _GEN_193; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_62 = _GEN_62[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_194 = {{61'd0}, mout_62}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2567 = _T_2566 + _GEN_194; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_63 = _GEN_63[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_195 = {{62'd0}, mout_63}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2568 = _T_2567 + _GEN_195; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_64 = _GEN_64[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_196 = {{63'd0}, mout_64}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2569 = _T_2568 + _GEN_196; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_65 = _GEN_65[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_197 = {{64'd0}, mout_65}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2570 = _T_2569 + _GEN_197; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_66 = _GEN_66[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_198 = {{65'd0}, mout_66}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2571 = _T_2570 + _GEN_198; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_67 = _GEN_67[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_199 = {{66'd0}, mout_67}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2572 = _T_2571 + _GEN_199; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_68 = _GEN_68[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_200 = {{67'd0}, mout_68}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2573 = _T_2572 + _GEN_200; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_69 = _GEN_69[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_201 = {{68'd0}, mout_69}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2574 = _T_2573 + _GEN_201; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_70 = _GEN_70[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_202 = {{69'd0}, mout_70}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2575 = _T_2574 + _GEN_202; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_71 = _GEN_71[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_203 = {{70'd0}, mout_71}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2576 = _T_2575 + _GEN_203; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_72 = _GEN_72[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_204 = {{71'd0}, mout_72}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2577 = _T_2576 + _GEN_204; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_73 = _GEN_73[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_205 = {{72'd0}, mout_73}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2578 = _T_2577 + _GEN_205; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_74 = _GEN_74[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_206 = {{73'd0}, mout_74}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2579 = _T_2578 + _GEN_206; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_75 = _GEN_75[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_207 = {{74'd0}, mout_75}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2580 = _T_2579 + _GEN_207; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_76 = _GEN_76[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_208 = {{75'd0}, mout_76}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2581 = _T_2580 + _GEN_208; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_77 = _GEN_77[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_209 = {{76'd0}, mout_77}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2582 = _T_2581 + _GEN_209; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_78 = _GEN_78[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_210 = {{77'd0}, mout_78}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2583 = _T_2582 + _GEN_210; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_79 = _GEN_79[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_211 = {{78'd0}, mout_79}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2584 = _T_2583 + _GEN_211; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_80 = _GEN_80[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_212 = {{79'd0}, mout_80}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2585 = _T_2584 + _GEN_212; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_81 = _GEN_81[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_213 = {{80'd0}, mout_81}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2586 = _T_2585 + _GEN_213; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_82 = _GEN_82[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_214 = {{81'd0}, mout_82}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2587 = _T_2586 + _GEN_214; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_83 = _GEN_83[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_215 = {{82'd0}, mout_83}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2588 = _T_2587 + _GEN_215; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_84 = _GEN_84[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_216 = {{83'd0}, mout_84}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2589 = _T_2588 + _GEN_216; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_85 = _GEN_85[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_217 = {{84'd0}, mout_85}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2590 = _T_2589 + _GEN_217; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_86 = _GEN_86[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_218 = {{85'd0}, mout_86}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2591 = _T_2590 + _GEN_218; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_87 = _GEN_87[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_219 = {{86'd0}, mout_87}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2592 = _T_2591 + _GEN_219; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_88 = _GEN_88[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_220 = {{87'd0}, mout_88}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2593 = _T_2592 + _GEN_220; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_89 = _GEN_89[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_221 = {{88'd0}, mout_89}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2594 = _T_2593 + _GEN_221; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_90 = _GEN_90[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_222 = {{89'd0}, mout_90}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2595 = _T_2594 + _GEN_222; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_91 = _GEN_91[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_223 = {{90'd0}, mout_91}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2596 = _T_2595 + _GEN_223; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_92 = _GEN_92[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_224 = {{91'd0}, mout_92}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2597 = _T_2596 + _GEN_224; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_93 = _GEN_93[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_225 = {{92'd0}, mout_93}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2598 = _T_2597 + _GEN_225; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_94 = _GEN_94[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_226 = {{93'd0}, mout_94}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2599 = _T_2598 + _GEN_226; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_95 = _GEN_95[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_227 = {{94'd0}, mout_95}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2600 = _T_2599 + _GEN_227; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_96 = _GEN_96[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_228 = {{95'd0}, mout_96}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2601 = _T_2600 + _GEN_228; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_97 = _GEN_97[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_229 = {{96'd0}, mout_97}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2602 = _T_2601 + _GEN_229; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_98 = _GEN_98[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_230 = {{97'd0}, mout_98}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2603 = _T_2602 + _GEN_230; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_99 = _GEN_99[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_231 = {{98'd0}, mout_99}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2604 = _T_2603 + _GEN_231; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_100 = _GEN_100[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_232 = {{99'd0}, mout_100}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2605 = _T_2604 + _GEN_232; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_101 = _GEN_101[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_233 = {{100'd0}, mout_101}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2606 = _T_2605 + _GEN_233; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_102 = _GEN_102[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_234 = {{101'd0}, mout_102}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2607 = _T_2606 + _GEN_234; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_103 = _GEN_103[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_235 = {{102'd0}, mout_103}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2608 = _T_2607 + _GEN_235; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_104 = _GEN_104[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_236 = {{103'd0}, mout_104}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2609 = _T_2608 + _GEN_236; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_105 = _GEN_105[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_237 = {{104'd0}, mout_105}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2610 = _T_2609 + _GEN_237; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_106 = _GEN_106[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_238 = {{105'd0}, mout_106}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2611 = _T_2610 + _GEN_238; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_107 = _GEN_107[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_239 = {{106'd0}, mout_107}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2612 = _T_2611 + _GEN_239; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_108 = _GEN_108[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_240 = {{107'd0}, mout_108}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2613 = _T_2612 + _GEN_240; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_109 = _GEN_109[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_241 = {{108'd0}, mout_109}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2614 = _T_2613 + _GEN_241; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_110 = _GEN_110[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_242 = {{109'd0}, mout_110}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2615 = _T_2614 + _GEN_242; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_111 = _GEN_111[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_243 = {{110'd0}, mout_111}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2616 = _T_2615 + _GEN_243; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_112 = _GEN_112[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_244 = {{111'd0}, mout_112}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2617 = _T_2616 + _GEN_244; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_113 = _GEN_113[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_245 = {{112'd0}, mout_113}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2618 = _T_2617 + _GEN_245; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_114 = _GEN_114[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_246 = {{113'd0}, mout_114}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2619 = _T_2618 + _GEN_246; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_115 = _GEN_115[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_247 = {{114'd0}, mout_115}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2620 = _T_2619 + _GEN_247; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_116 = _GEN_116[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_248 = {{115'd0}, mout_116}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2621 = _T_2620 + _GEN_248; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_117 = _GEN_117[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_249 = {{116'd0}, mout_117}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2622 = _T_2621 + _GEN_249; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_118 = _GEN_118[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_250 = {{117'd0}, mout_118}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2623 = _T_2622 + _GEN_250; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_119 = _GEN_119[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_251 = {{118'd0}, mout_119}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2624 = _T_2623 + _GEN_251; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_120 = _GEN_120[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_252 = {{119'd0}, mout_120}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2625 = _T_2624 + _GEN_252; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_121 = _GEN_121[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_253 = {{120'd0}, mout_121}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2626 = _T_2625 + _GEN_253; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_122 = _GEN_122[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_254 = {{121'd0}, mout_122}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2627 = _T_2626 + _GEN_254; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_123 = _GEN_123[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_255 = {{122'd0}, mout_123}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2628 = _T_2627 + _GEN_255; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_124 = _GEN_124[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_256 = {{123'd0}, mout_124}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2629 = _T_2628 + _GEN_256; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_125 = _GEN_125[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_257 = {{124'd0}, mout_125}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2630 = _T_2629 + _GEN_257; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_126 = _GEN_126[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_258 = {{125'd0}, mout_126}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign _T_2631 = _T_2630 + _GEN_258; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign mout_127 = _GEN_127[15:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 48:23 NV_NVDLA_CMAC_CORE_mac.scala 52:22 NV_NVDLA_CMAC_CORE_mac.scala 55:22]
  assign _GEN_259 = {{126'd0}, mout_127}; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign sum_out = _T_2631 + _GEN_259; // @[NV_NVDLA_CMAC_CORE_mac.scala 59:32]
  assign pp_pvld_d0 = io_dat_actv_pvld_0 & io_wt_actv_pvld_0; // @[NV_NVDLA_CMAC_CORE_mac.scala 62:41]
  assign io_mac_out_data = _T_2637[22:0]; // @[NV_NVDLA_CMAC_CORE_mac.scala 64:21]
  assign io_mac_out_pvld = _T_2643; // @[NV_NVDLA_CMAC_CORE_mac.scala 65:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  _T_2633 = _RAND_0[142:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {5{`RANDOM}};
  _T_2635 = _RAND_1[142:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {5{`RANDOM}};
  _T_2637 = _RAND_2[142:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2639 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2641 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2643 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (pp_pvld_d0) begin
      _T_2633 <= sum_out;
    end
    if (pp_pvld_d0) begin
      _T_2635 <= _T_2633;
    end
    if (pp_pvld_d0) begin
      _T_2637 <= _T_2635;
    end
    if (pp_pvld_d0) begin
      _T_2639 <= pp_pvld_d0;
    end
    if (pp_pvld_d0) begin
      _T_2641 <= _T_2639;
    end
    if (pp_pvld_d0) begin
      _T_2643 <= _T_2641;
    end
  end
endmodule
module NV_NVDLA_CMAC_CORE_rt_out(
  input         clock,
  input         reset,
  input  [22:0] io_out_data_0,
  input         io_out_mask_0,
  input  [8:0]  io_out_pd,
  input         io_out_pvld,
  output [22:0] io_mac2accu_data_0,
  output        io_mac2accu_mask_0,
  output [8:0]  io_mac2accu_pd,
  output        io_mac2accu_pvld,
  output        io_dp2reg_done
);
  reg  out_rt_pvld_d_1; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 50:67]
  reg [31:0] _RAND_0;
  reg  out_rt_pvld_d_2; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 50:67]
  reg [31:0] _RAND_1;
  reg  out_rt_mask_d_1_0; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 53:67]
  reg [31:0] _RAND_2;
  reg  out_rt_mask_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 53:67]
  reg [31:0] _RAND_3;
  reg [8:0] out_rt_pd_d_1; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 56:65]
  reg [31:0] _RAND_4;
  reg [8:0] out_rt_pd_d_2; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 56:65]
  reg [31:0] _RAND_5;
  reg [22:0] out_rt_data_d_1_0; // @[retiming.scala 9:92]
  reg [31:0] _RAND_6;
  reg [22:0] out_rt_data_d_2_0; // @[retiming.scala 9:92]
  reg [31:0] _RAND_7;
  reg  dp2reg_done_d_1; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 61:67]
  reg [31:0] _RAND_8;
  reg  dp2reg_done_d_2; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 61:67]
  reg [31:0] _RAND_9;
  wire  _T_138; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 68:34]
  wire  _T_139; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 68:88]
  wire  _T_140; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 68:78]
  wire  dp2reg_done_d_0; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 68:133]
  wire [8:0] _GEN_0; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 75:31]
  wire [8:0] _GEN_2; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 75:31]
  assign _T_138 = io_out_pd[8]; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 68:34]
  assign _T_139 = io_out_pd[6]; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 68:88]
  assign _T_140 = _T_138 & _T_139; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 68:78]
  assign dp2reg_done_d_0 = _T_140 & io_out_pvld; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 68:133]
  assign _GEN_0 = io_out_pvld ? io_out_pd : out_rt_pd_d_1; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 75:31]
  assign _GEN_2 = out_rt_pvld_d_1 ? out_rt_pd_d_1 : out_rt_pd_d_2; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 75:31]
  assign io_mac2accu_data_0 = out_rt_data_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 89:22]
  assign io_mac2accu_mask_0 = out_rt_mask_d_2_0; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 87:22]
  assign io_mac2accu_pd = out_rt_pd_d_2; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 88:20]
  assign io_mac2accu_pvld = out_rt_pvld_d_2; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 86:22]
  assign io_dp2reg_done = dp2reg_done_d_2; // @[NV_NVDLA_CMAC_CORE_rt_out.scala 91:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_rt_pvld_d_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_rt_pvld_d_2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_rt_mask_d_1_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_rt_mask_d_2_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_rt_pd_d_1 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_rt_pd_d_2 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_rt_data_d_1_0 = _RAND_6[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_rt_data_d_2_0 = _RAND_7[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  dp2reg_done_d_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  dp2reg_done_d_2 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_rt_pvld_d_1 <= 1'h0;
    end else begin
      out_rt_pvld_d_1 <= io_out_pvld;
    end
    if (reset) begin
      out_rt_pvld_d_2 <= 1'h0;
    end else begin
      out_rt_pvld_d_2 <= out_rt_pvld_d_1;
    end
    if (reset) begin
      out_rt_mask_d_1_0 <= 1'h0;
    end else begin
      out_rt_mask_d_1_0 <= io_out_mask_0;
    end
    if (reset) begin
      out_rt_mask_d_2_0 <= 1'h0;
    end else begin
      out_rt_mask_d_2_0 <= out_rt_mask_d_1_0;
    end
    if (reset) begin
      out_rt_pd_d_1 <= 9'h0;
    end else begin
      if (io_out_pvld) begin
        out_rt_pd_d_1 <= io_out_pd;
      end
    end
    if (reset) begin
      out_rt_pd_d_2 <= 9'h0;
    end else begin
      if (out_rt_pvld_d_1) begin
        out_rt_pd_d_2 <= out_rt_pd_d_1;
      end
    end
    if (io_out_mask_0) begin
      out_rt_data_d_1_0 <= io_out_data_0;
    end
    if (out_rt_mask_d_1_0) begin
      out_rt_data_d_2_0 <= out_rt_data_d_1_0;
    end
    if (reset) begin
      dp2reg_done_d_1 <= 1'h0;
    end else begin
      dp2reg_done_d_1 <= dp2reg_done_d_0;
    end
    if (reset) begin
      dp2reg_done_d_2 <= 1'h0;
    end else begin
      dp2reg_done_d_2 <= dp2reg_done_d_1;
    end
  end
endmodule
module NV_NVDLA_CMAC_core(
  input         clock,
  input         reset,
  input         io_sc2mac_dat_pvld,
  input         io_sc2mac_dat_mask_0,
  input         io_sc2mac_dat_mask_1,
  input         io_sc2mac_dat_mask_2,
  input         io_sc2mac_dat_mask_3,
  input         io_sc2mac_dat_mask_4,
  input         io_sc2mac_dat_mask_5,
  input         io_sc2mac_dat_mask_6,
  input         io_sc2mac_dat_mask_7,
  input         io_sc2mac_dat_mask_8,
  input         io_sc2mac_dat_mask_9,
  input         io_sc2mac_dat_mask_10,
  input         io_sc2mac_dat_mask_11,
  input         io_sc2mac_dat_mask_12,
  input         io_sc2mac_dat_mask_13,
  input         io_sc2mac_dat_mask_14,
  input         io_sc2mac_dat_mask_15,
  input         io_sc2mac_dat_mask_16,
  input         io_sc2mac_dat_mask_17,
  input         io_sc2mac_dat_mask_18,
  input         io_sc2mac_dat_mask_19,
  input         io_sc2mac_dat_mask_20,
  input         io_sc2mac_dat_mask_21,
  input         io_sc2mac_dat_mask_22,
  input         io_sc2mac_dat_mask_23,
  input         io_sc2mac_dat_mask_24,
  input         io_sc2mac_dat_mask_25,
  input         io_sc2mac_dat_mask_26,
  input         io_sc2mac_dat_mask_27,
  input         io_sc2mac_dat_mask_28,
  input         io_sc2mac_dat_mask_29,
  input         io_sc2mac_dat_mask_30,
  input         io_sc2mac_dat_mask_31,
  input         io_sc2mac_dat_mask_32,
  input         io_sc2mac_dat_mask_33,
  input         io_sc2mac_dat_mask_34,
  input         io_sc2mac_dat_mask_35,
  input         io_sc2mac_dat_mask_36,
  input         io_sc2mac_dat_mask_37,
  input         io_sc2mac_dat_mask_38,
  input         io_sc2mac_dat_mask_39,
  input         io_sc2mac_dat_mask_40,
  input         io_sc2mac_dat_mask_41,
  input         io_sc2mac_dat_mask_42,
  input         io_sc2mac_dat_mask_43,
  input         io_sc2mac_dat_mask_44,
  input         io_sc2mac_dat_mask_45,
  input         io_sc2mac_dat_mask_46,
  input         io_sc2mac_dat_mask_47,
  input         io_sc2mac_dat_mask_48,
  input         io_sc2mac_dat_mask_49,
  input         io_sc2mac_dat_mask_50,
  input         io_sc2mac_dat_mask_51,
  input         io_sc2mac_dat_mask_52,
  input         io_sc2mac_dat_mask_53,
  input         io_sc2mac_dat_mask_54,
  input         io_sc2mac_dat_mask_55,
  input         io_sc2mac_dat_mask_56,
  input         io_sc2mac_dat_mask_57,
  input         io_sc2mac_dat_mask_58,
  input         io_sc2mac_dat_mask_59,
  input         io_sc2mac_dat_mask_60,
  input         io_sc2mac_dat_mask_61,
  input         io_sc2mac_dat_mask_62,
  input         io_sc2mac_dat_mask_63,
  input         io_sc2mac_dat_mask_64,
  input         io_sc2mac_dat_mask_65,
  input         io_sc2mac_dat_mask_66,
  input         io_sc2mac_dat_mask_67,
  input         io_sc2mac_dat_mask_68,
  input         io_sc2mac_dat_mask_69,
  input         io_sc2mac_dat_mask_70,
  input         io_sc2mac_dat_mask_71,
  input         io_sc2mac_dat_mask_72,
  input         io_sc2mac_dat_mask_73,
  input         io_sc2mac_dat_mask_74,
  input         io_sc2mac_dat_mask_75,
  input         io_sc2mac_dat_mask_76,
  input         io_sc2mac_dat_mask_77,
  input         io_sc2mac_dat_mask_78,
  input         io_sc2mac_dat_mask_79,
  input         io_sc2mac_dat_mask_80,
  input         io_sc2mac_dat_mask_81,
  input         io_sc2mac_dat_mask_82,
  input         io_sc2mac_dat_mask_83,
  input         io_sc2mac_dat_mask_84,
  input         io_sc2mac_dat_mask_85,
  input         io_sc2mac_dat_mask_86,
  input         io_sc2mac_dat_mask_87,
  input         io_sc2mac_dat_mask_88,
  input         io_sc2mac_dat_mask_89,
  input         io_sc2mac_dat_mask_90,
  input         io_sc2mac_dat_mask_91,
  input         io_sc2mac_dat_mask_92,
  input         io_sc2mac_dat_mask_93,
  input         io_sc2mac_dat_mask_94,
  input         io_sc2mac_dat_mask_95,
  input         io_sc2mac_dat_mask_96,
  input         io_sc2mac_dat_mask_97,
  input         io_sc2mac_dat_mask_98,
  input         io_sc2mac_dat_mask_99,
  input         io_sc2mac_dat_mask_100,
  input         io_sc2mac_dat_mask_101,
  input         io_sc2mac_dat_mask_102,
  input         io_sc2mac_dat_mask_103,
  input         io_sc2mac_dat_mask_104,
  input         io_sc2mac_dat_mask_105,
  input         io_sc2mac_dat_mask_106,
  input         io_sc2mac_dat_mask_107,
  input         io_sc2mac_dat_mask_108,
  input         io_sc2mac_dat_mask_109,
  input         io_sc2mac_dat_mask_110,
  input         io_sc2mac_dat_mask_111,
  input         io_sc2mac_dat_mask_112,
  input         io_sc2mac_dat_mask_113,
  input         io_sc2mac_dat_mask_114,
  input         io_sc2mac_dat_mask_115,
  input         io_sc2mac_dat_mask_116,
  input         io_sc2mac_dat_mask_117,
  input         io_sc2mac_dat_mask_118,
  input         io_sc2mac_dat_mask_119,
  input         io_sc2mac_dat_mask_120,
  input         io_sc2mac_dat_mask_121,
  input         io_sc2mac_dat_mask_122,
  input         io_sc2mac_dat_mask_123,
  input         io_sc2mac_dat_mask_124,
  input         io_sc2mac_dat_mask_125,
  input         io_sc2mac_dat_mask_126,
  input         io_sc2mac_dat_mask_127,
  input  [7:0]  io_sc2mac_dat_data_0,
  input  [7:0]  io_sc2mac_dat_data_1,
  input  [7:0]  io_sc2mac_dat_data_2,
  input  [7:0]  io_sc2mac_dat_data_3,
  input  [7:0]  io_sc2mac_dat_data_4,
  input  [7:0]  io_sc2mac_dat_data_5,
  input  [7:0]  io_sc2mac_dat_data_6,
  input  [7:0]  io_sc2mac_dat_data_7,
  input  [7:0]  io_sc2mac_dat_data_8,
  input  [7:0]  io_sc2mac_dat_data_9,
  input  [7:0]  io_sc2mac_dat_data_10,
  input  [7:0]  io_sc2mac_dat_data_11,
  input  [7:0]  io_sc2mac_dat_data_12,
  input  [7:0]  io_sc2mac_dat_data_13,
  input  [7:0]  io_sc2mac_dat_data_14,
  input  [7:0]  io_sc2mac_dat_data_15,
  input  [7:0]  io_sc2mac_dat_data_16,
  input  [7:0]  io_sc2mac_dat_data_17,
  input  [7:0]  io_sc2mac_dat_data_18,
  input  [7:0]  io_sc2mac_dat_data_19,
  input  [7:0]  io_sc2mac_dat_data_20,
  input  [7:0]  io_sc2mac_dat_data_21,
  input  [7:0]  io_sc2mac_dat_data_22,
  input  [7:0]  io_sc2mac_dat_data_23,
  input  [7:0]  io_sc2mac_dat_data_24,
  input  [7:0]  io_sc2mac_dat_data_25,
  input  [7:0]  io_sc2mac_dat_data_26,
  input  [7:0]  io_sc2mac_dat_data_27,
  input  [7:0]  io_sc2mac_dat_data_28,
  input  [7:0]  io_sc2mac_dat_data_29,
  input  [7:0]  io_sc2mac_dat_data_30,
  input  [7:0]  io_sc2mac_dat_data_31,
  input  [7:0]  io_sc2mac_dat_data_32,
  input  [7:0]  io_sc2mac_dat_data_33,
  input  [7:0]  io_sc2mac_dat_data_34,
  input  [7:0]  io_sc2mac_dat_data_35,
  input  [7:0]  io_sc2mac_dat_data_36,
  input  [7:0]  io_sc2mac_dat_data_37,
  input  [7:0]  io_sc2mac_dat_data_38,
  input  [7:0]  io_sc2mac_dat_data_39,
  input  [7:0]  io_sc2mac_dat_data_40,
  input  [7:0]  io_sc2mac_dat_data_41,
  input  [7:0]  io_sc2mac_dat_data_42,
  input  [7:0]  io_sc2mac_dat_data_43,
  input  [7:0]  io_sc2mac_dat_data_44,
  input  [7:0]  io_sc2mac_dat_data_45,
  input  [7:0]  io_sc2mac_dat_data_46,
  input  [7:0]  io_sc2mac_dat_data_47,
  input  [7:0]  io_sc2mac_dat_data_48,
  input  [7:0]  io_sc2mac_dat_data_49,
  input  [7:0]  io_sc2mac_dat_data_50,
  input  [7:0]  io_sc2mac_dat_data_51,
  input  [7:0]  io_sc2mac_dat_data_52,
  input  [7:0]  io_sc2mac_dat_data_53,
  input  [7:0]  io_sc2mac_dat_data_54,
  input  [7:0]  io_sc2mac_dat_data_55,
  input  [7:0]  io_sc2mac_dat_data_56,
  input  [7:0]  io_sc2mac_dat_data_57,
  input  [7:0]  io_sc2mac_dat_data_58,
  input  [7:0]  io_sc2mac_dat_data_59,
  input  [7:0]  io_sc2mac_dat_data_60,
  input  [7:0]  io_sc2mac_dat_data_61,
  input  [7:0]  io_sc2mac_dat_data_62,
  input  [7:0]  io_sc2mac_dat_data_63,
  input  [7:0]  io_sc2mac_dat_data_64,
  input  [7:0]  io_sc2mac_dat_data_65,
  input  [7:0]  io_sc2mac_dat_data_66,
  input  [7:0]  io_sc2mac_dat_data_67,
  input  [7:0]  io_sc2mac_dat_data_68,
  input  [7:0]  io_sc2mac_dat_data_69,
  input  [7:0]  io_sc2mac_dat_data_70,
  input  [7:0]  io_sc2mac_dat_data_71,
  input  [7:0]  io_sc2mac_dat_data_72,
  input  [7:0]  io_sc2mac_dat_data_73,
  input  [7:0]  io_sc2mac_dat_data_74,
  input  [7:0]  io_sc2mac_dat_data_75,
  input  [7:0]  io_sc2mac_dat_data_76,
  input  [7:0]  io_sc2mac_dat_data_77,
  input  [7:0]  io_sc2mac_dat_data_78,
  input  [7:0]  io_sc2mac_dat_data_79,
  input  [7:0]  io_sc2mac_dat_data_80,
  input  [7:0]  io_sc2mac_dat_data_81,
  input  [7:0]  io_sc2mac_dat_data_82,
  input  [7:0]  io_sc2mac_dat_data_83,
  input  [7:0]  io_sc2mac_dat_data_84,
  input  [7:0]  io_sc2mac_dat_data_85,
  input  [7:0]  io_sc2mac_dat_data_86,
  input  [7:0]  io_sc2mac_dat_data_87,
  input  [7:0]  io_sc2mac_dat_data_88,
  input  [7:0]  io_sc2mac_dat_data_89,
  input  [7:0]  io_sc2mac_dat_data_90,
  input  [7:0]  io_sc2mac_dat_data_91,
  input  [7:0]  io_sc2mac_dat_data_92,
  input  [7:0]  io_sc2mac_dat_data_93,
  input  [7:0]  io_sc2mac_dat_data_94,
  input  [7:0]  io_sc2mac_dat_data_95,
  input  [7:0]  io_sc2mac_dat_data_96,
  input  [7:0]  io_sc2mac_dat_data_97,
  input  [7:0]  io_sc2mac_dat_data_98,
  input  [7:0]  io_sc2mac_dat_data_99,
  input  [7:0]  io_sc2mac_dat_data_100,
  input  [7:0]  io_sc2mac_dat_data_101,
  input  [7:0]  io_sc2mac_dat_data_102,
  input  [7:0]  io_sc2mac_dat_data_103,
  input  [7:0]  io_sc2mac_dat_data_104,
  input  [7:0]  io_sc2mac_dat_data_105,
  input  [7:0]  io_sc2mac_dat_data_106,
  input  [7:0]  io_sc2mac_dat_data_107,
  input  [7:0]  io_sc2mac_dat_data_108,
  input  [7:0]  io_sc2mac_dat_data_109,
  input  [7:0]  io_sc2mac_dat_data_110,
  input  [7:0]  io_sc2mac_dat_data_111,
  input  [7:0]  io_sc2mac_dat_data_112,
  input  [7:0]  io_sc2mac_dat_data_113,
  input  [7:0]  io_sc2mac_dat_data_114,
  input  [7:0]  io_sc2mac_dat_data_115,
  input  [7:0]  io_sc2mac_dat_data_116,
  input  [7:0]  io_sc2mac_dat_data_117,
  input  [7:0]  io_sc2mac_dat_data_118,
  input  [7:0]  io_sc2mac_dat_data_119,
  input  [7:0]  io_sc2mac_dat_data_120,
  input  [7:0]  io_sc2mac_dat_data_121,
  input  [7:0]  io_sc2mac_dat_data_122,
  input  [7:0]  io_sc2mac_dat_data_123,
  input  [7:0]  io_sc2mac_dat_data_124,
  input  [7:0]  io_sc2mac_dat_data_125,
  input  [7:0]  io_sc2mac_dat_data_126,
  input  [7:0]  io_sc2mac_dat_data_127,
  input  [8:0]  io_sc2mac_dat_pd,
  input         io_sc2mac_wt_pvld,
  input         io_sc2mac_wt_mask_0,
  input         io_sc2mac_wt_mask_1,
  input         io_sc2mac_wt_mask_2,
  input         io_sc2mac_wt_mask_3,
  input         io_sc2mac_wt_mask_4,
  input         io_sc2mac_wt_mask_5,
  input         io_sc2mac_wt_mask_6,
  input         io_sc2mac_wt_mask_7,
  input         io_sc2mac_wt_mask_8,
  input         io_sc2mac_wt_mask_9,
  input         io_sc2mac_wt_mask_10,
  input         io_sc2mac_wt_mask_11,
  input         io_sc2mac_wt_mask_12,
  input         io_sc2mac_wt_mask_13,
  input         io_sc2mac_wt_mask_14,
  input         io_sc2mac_wt_mask_15,
  input         io_sc2mac_wt_mask_16,
  input         io_sc2mac_wt_mask_17,
  input         io_sc2mac_wt_mask_18,
  input         io_sc2mac_wt_mask_19,
  input         io_sc2mac_wt_mask_20,
  input         io_sc2mac_wt_mask_21,
  input         io_sc2mac_wt_mask_22,
  input         io_sc2mac_wt_mask_23,
  input         io_sc2mac_wt_mask_24,
  input         io_sc2mac_wt_mask_25,
  input         io_sc2mac_wt_mask_26,
  input         io_sc2mac_wt_mask_27,
  input         io_sc2mac_wt_mask_28,
  input         io_sc2mac_wt_mask_29,
  input         io_sc2mac_wt_mask_30,
  input         io_sc2mac_wt_mask_31,
  input         io_sc2mac_wt_mask_32,
  input         io_sc2mac_wt_mask_33,
  input         io_sc2mac_wt_mask_34,
  input         io_sc2mac_wt_mask_35,
  input         io_sc2mac_wt_mask_36,
  input         io_sc2mac_wt_mask_37,
  input         io_sc2mac_wt_mask_38,
  input         io_sc2mac_wt_mask_39,
  input         io_sc2mac_wt_mask_40,
  input         io_sc2mac_wt_mask_41,
  input         io_sc2mac_wt_mask_42,
  input         io_sc2mac_wt_mask_43,
  input         io_sc2mac_wt_mask_44,
  input         io_sc2mac_wt_mask_45,
  input         io_sc2mac_wt_mask_46,
  input         io_sc2mac_wt_mask_47,
  input         io_sc2mac_wt_mask_48,
  input         io_sc2mac_wt_mask_49,
  input         io_sc2mac_wt_mask_50,
  input         io_sc2mac_wt_mask_51,
  input         io_sc2mac_wt_mask_52,
  input         io_sc2mac_wt_mask_53,
  input         io_sc2mac_wt_mask_54,
  input         io_sc2mac_wt_mask_55,
  input         io_sc2mac_wt_mask_56,
  input         io_sc2mac_wt_mask_57,
  input         io_sc2mac_wt_mask_58,
  input         io_sc2mac_wt_mask_59,
  input         io_sc2mac_wt_mask_60,
  input         io_sc2mac_wt_mask_61,
  input         io_sc2mac_wt_mask_62,
  input         io_sc2mac_wt_mask_63,
  input         io_sc2mac_wt_mask_64,
  input         io_sc2mac_wt_mask_65,
  input         io_sc2mac_wt_mask_66,
  input         io_sc2mac_wt_mask_67,
  input         io_sc2mac_wt_mask_68,
  input         io_sc2mac_wt_mask_69,
  input         io_sc2mac_wt_mask_70,
  input         io_sc2mac_wt_mask_71,
  input         io_sc2mac_wt_mask_72,
  input         io_sc2mac_wt_mask_73,
  input         io_sc2mac_wt_mask_74,
  input         io_sc2mac_wt_mask_75,
  input         io_sc2mac_wt_mask_76,
  input         io_sc2mac_wt_mask_77,
  input         io_sc2mac_wt_mask_78,
  input         io_sc2mac_wt_mask_79,
  input         io_sc2mac_wt_mask_80,
  input         io_sc2mac_wt_mask_81,
  input         io_sc2mac_wt_mask_82,
  input         io_sc2mac_wt_mask_83,
  input         io_sc2mac_wt_mask_84,
  input         io_sc2mac_wt_mask_85,
  input         io_sc2mac_wt_mask_86,
  input         io_sc2mac_wt_mask_87,
  input         io_sc2mac_wt_mask_88,
  input         io_sc2mac_wt_mask_89,
  input         io_sc2mac_wt_mask_90,
  input         io_sc2mac_wt_mask_91,
  input         io_sc2mac_wt_mask_92,
  input         io_sc2mac_wt_mask_93,
  input         io_sc2mac_wt_mask_94,
  input         io_sc2mac_wt_mask_95,
  input         io_sc2mac_wt_mask_96,
  input         io_sc2mac_wt_mask_97,
  input         io_sc2mac_wt_mask_98,
  input         io_sc2mac_wt_mask_99,
  input         io_sc2mac_wt_mask_100,
  input         io_sc2mac_wt_mask_101,
  input         io_sc2mac_wt_mask_102,
  input         io_sc2mac_wt_mask_103,
  input         io_sc2mac_wt_mask_104,
  input         io_sc2mac_wt_mask_105,
  input         io_sc2mac_wt_mask_106,
  input         io_sc2mac_wt_mask_107,
  input         io_sc2mac_wt_mask_108,
  input         io_sc2mac_wt_mask_109,
  input         io_sc2mac_wt_mask_110,
  input         io_sc2mac_wt_mask_111,
  input         io_sc2mac_wt_mask_112,
  input         io_sc2mac_wt_mask_113,
  input         io_sc2mac_wt_mask_114,
  input         io_sc2mac_wt_mask_115,
  input         io_sc2mac_wt_mask_116,
  input         io_sc2mac_wt_mask_117,
  input         io_sc2mac_wt_mask_118,
  input         io_sc2mac_wt_mask_119,
  input         io_sc2mac_wt_mask_120,
  input         io_sc2mac_wt_mask_121,
  input         io_sc2mac_wt_mask_122,
  input         io_sc2mac_wt_mask_123,
  input         io_sc2mac_wt_mask_124,
  input         io_sc2mac_wt_mask_125,
  input         io_sc2mac_wt_mask_126,
  input         io_sc2mac_wt_mask_127,
  input  [7:0]  io_sc2mac_wt_data_0,
  input  [7:0]  io_sc2mac_wt_data_1,
  input  [7:0]  io_sc2mac_wt_data_2,
  input  [7:0]  io_sc2mac_wt_data_3,
  input  [7:0]  io_sc2mac_wt_data_4,
  input  [7:0]  io_sc2mac_wt_data_5,
  input  [7:0]  io_sc2mac_wt_data_6,
  input  [7:0]  io_sc2mac_wt_data_7,
  input  [7:0]  io_sc2mac_wt_data_8,
  input  [7:0]  io_sc2mac_wt_data_9,
  input  [7:0]  io_sc2mac_wt_data_10,
  input  [7:0]  io_sc2mac_wt_data_11,
  input  [7:0]  io_sc2mac_wt_data_12,
  input  [7:0]  io_sc2mac_wt_data_13,
  input  [7:0]  io_sc2mac_wt_data_14,
  input  [7:0]  io_sc2mac_wt_data_15,
  input  [7:0]  io_sc2mac_wt_data_16,
  input  [7:0]  io_sc2mac_wt_data_17,
  input  [7:0]  io_sc2mac_wt_data_18,
  input  [7:0]  io_sc2mac_wt_data_19,
  input  [7:0]  io_sc2mac_wt_data_20,
  input  [7:0]  io_sc2mac_wt_data_21,
  input  [7:0]  io_sc2mac_wt_data_22,
  input  [7:0]  io_sc2mac_wt_data_23,
  input  [7:0]  io_sc2mac_wt_data_24,
  input  [7:0]  io_sc2mac_wt_data_25,
  input  [7:0]  io_sc2mac_wt_data_26,
  input  [7:0]  io_sc2mac_wt_data_27,
  input  [7:0]  io_sc2mac_wt_data_28,
  input  [7:0]  io_sc2mac_wt_data_29,
  input  [7:0]  io_sc2mac_wt_data_30,
  input  [7:0]  io_sc2mac_wt_data_31,
  input  [7:0]  io_sc2mac_wt_data_32,
  input  [7:0]  io_sc2mac_wt_data_33,
  input  [7:0]  io_sc2mac_wt_data_34,
  input  [7:0]  io_sc2mac_wt_data_35,
  input  [7:0]  io_sc2mac_wt_data_36,
  input  [7:0]  io_sc2mac_wt_data_37,
  input  [7:0]  io_sc2mac_wt_data_38,
  input  [7:0]  io_sc2mac_wt_data_39,
  input  [7:0]  io_sc2mac_wt_data_40,
  input  [7:0]  io_sc2mac_wt_data_41,
  input  [7:0]  io_sc2mac_wt_data_42,
  input  [7:0]  io_sc2mac_wt_data_43,
  input  [7:0]  io_sc2mac_wt_data_44,
  input  [7:0]  io_sc2mac_wt_data_45,
  input  [7:0]  io_sc2mac_wt_data_46,
  input  [7:0]  io_sc2mac_wt_data_47,
  input  [7:0]  io_sc2mac_wt_data_48,
  input  [7:0]  io_sc2mac_wt_data_49,
  input  [7:0]  io_sc2mac_wt_data_50,
  input  [7:0]  io_sc2mac_wt_data_51,
  input  [7:0]  io_sc2mac_wt_data_52,
  input  [7:0]  io_sc2mac_wt_data_53,
  input  [7:0]  io_sc2mac_wt_data_54,
  input  [7:0]  io_sc2mac_wt_data_55,
  input  [7:0]  io_sc2mac_wt_data_56,
  input  [7:0]  io_sc2mac_wt_data_57,
  input  [7:0]  io_sc2mac_wt_data_58,
  input  [7:0]  io_sc2mac_wt_data_59,
  input  [7:0]  io_sc2mac_wt_data_60,
  input  [7:0]  io_sc2mac_wt_data_61,
  input  [7:0]  io_sc2mac_wt_data_62,
  input  [7:0]  io_sc2mac_wt_data_63,
  input  [7:0]  io_sc2mac_wt_data_64,
  input  [7:0]  io_sc2mac_wt_data_65,
  input  [7:0]  io_sc2mac_wt_data_66,
  input  [7:0]  io_sc2mac_wt_data_67,
  input  [7:0]  io_sc2mac_wt_data_68,
  input  [7:0]  io_sc2mac_wt_data_69,
  input  [7:0]  io_sc2mac_wt_data_70,
  input  [7:0]  io_sc2mac_wt_data_71,
  input  [7:0]  io_sc2mac_wt_data_72,
  input  [7:0]  io_sc2mac_wt_data_73,
  input  [7:0]  io_sc2mac_wt_data_74,
  input  [7:0]  io_sc2mac_wt_data_75,
  input  [7:0]  io_sc2mac_wt_data_76,
  input  [7:0]  io_sc2mac_wt_data_77,
  input  [7:0]  io_sc2mac_wt_data_78,
  input  [7:0]  io_sc2mac_wt_data_79,
  input  [7:0]  io_sc2mac_wt_data_80,
  input  [7:0]  io_sc2mac_wt_data_81,
  input  [7:0]  io_sc2mac_wt_data_82,
  input  [7:0]  io_sc2mac_wt_data_83,
  input  [7:0]  io_sc2mac_wt_data_84,
  input  [7:0]  io_sc2mac_wt_data_85,
  input  [7:0]  io_sc2mac_wt_data_86,
  input  [7:0]  io_sc2mac_wt_data_87,
  input  [7:0]  io_sc2mac_wt_data_88,
  input  [7:0]  io_sc2mac_wt_data_89,
  input  [7:0]  io_sc2mac_wt_data_90,
  input  [7:0]  io_sc2mac_wt_data_91,
  input  [7:0]  io_sc2mac_wt_data_92,
  input  [7:0]  io_sc2mac_wt_data_93,
  input  [7:0]  io_sc2mac_wt_data_94,
  input  [7:0]  io_sc2mac_wt_data_95,
  input  [7:0]  io_sc2mac_wt_data_96,
  input  [7:0]  io_sc2mac_wt_data_97,
  input  [7:0]  io_sc2mac_wt_data_98,
  input  [7:0]  io_sc2mac_wt_data_99,
  input  [7:0]  io_sc2mac_wt_data_100,
  input  [7:0]  io_sc2mac_wt_data_101,
  input  [7:0]  io_sc2mac_wt_data_102,
  input  [7:0]  io_sc2mac_wt_data_103,
  input  [7:0]  io_sc2mac_wt_data_104,
  input  [7:0]  io_sc2mac_wt_data_105,
  input  [7:0]  io_sc2mac_wt_data_106,
  input  [7:0]  io_sc2mac_wt_data_107,
  input  [7:0]  io_sc2mac_wt_data_108,
  input  [7:0]  io_sc2mac_wt_data_109,
  input  [7:0]  io_sc2mac_wt_data_110,
  input  [7:0]  io_sc2mac_wt_data_111,
  input  [7:0]  io_sc2mac_wt_data_112,
  input  [7:0]  io_sc2mac_wt_data_113,
  input  [7:0]  io_sc2mac_wt_data_114,
  input  [7:0]  io_sc2mac_wt_data_115,
  input  [7:0]  io_sc2mac_wt_data_116,
  input  [7:0]  io_sc2mac_wt_data_117,
  input  [7:0]  io_sc2mac_wt_data_118,
  input  [7:0]  io_sc2mac_wt_data_119,
  input  [7:0]  io_sc2mac_wt_data_120,
  input  [7:0]  io_sc2mac_wt_data_121,
  input  [7:0]  io_sc2mac_wt_data_122,
  input  [7:0]  io_sc2mac_wt_data_123,
  input  [7:0]  io_sc2mac_wt_data_124,
  input  [7:0]  io_sc2mac_wt_data_125,
  input  [7:0]  io_sc2mac_wt_data_126,
  input  [7:0]  io_sc2mac_wt_data_127,
  input         io_sc2mac_wt_sel_0,
  output        io_mac2accu_pvld,
  output        io_mac2accu_mask_0,
  output [22:0] io_mac2accu_data_0,
  output [8:0]  io_mac2accu_pd,
  output        io_dp2reg_done
);
  wire  u_rt_in_clock; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_reset; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_1; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_2; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_3; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_4; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_5; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_6; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_7; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_8; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_9; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_10; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_11; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_12; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_13; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_14; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_15; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_16; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_17; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_18; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_19; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_20; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_21; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_22; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_23; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_24; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_25; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_26; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_27; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_28; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_29; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_30; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_31; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_32; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_33; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_34; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_35; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_36; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_37; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_38; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_39; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_40; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_41; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_42; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_43; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_44; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_45; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_46; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_47; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_48; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_49; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_50; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_51; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_52; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_53; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_54; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_55; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_56; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_57; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_58; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_59; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_60; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_61; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_62; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_63; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_64; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_65; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_66; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_67; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_68; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_69; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_70; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_71; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_72; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_73; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_74; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_75; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_76; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_77; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_78; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_79; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_80; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_81; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_82; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_83; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_84; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_85; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_86; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_87; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_88; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_89; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_90; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_91; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_92; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_93; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_94; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_95; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_96; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_97; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_98; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_99; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_100; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_101; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_102; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_103; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_104; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_105; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_106; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_107; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_108; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_109; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_110; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_111; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_112; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_113; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_114; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_115; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_116; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_117; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_118; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_119; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_120; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_121; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_122; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_123; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_124; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_125; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_126; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_dat_data_127; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_1; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_2; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_3; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_4; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_5; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_6; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_7; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_8; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_9; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_10; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_11; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_12; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_13; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_14; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_15; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_16; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_17; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_18; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_19; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_20; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_21; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_22; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_23; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_24; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_25; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_26; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_27; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_28; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_29; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_30; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_31; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_32; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_33; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_34; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_35; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_36; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_37; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_38; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_39; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_40; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_41; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_42; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_43; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_44; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_45; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_46; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_47; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_48; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_49; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_50; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_51; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_52; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_53; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_54; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_55; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_56; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_57; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_58; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_59; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_60; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_61; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_62; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_63; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_64; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_65; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_66; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_67; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_68; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_69; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_70; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_71; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_72; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_73; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_74; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_75; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_76; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_77; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_78; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_79; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_80; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_81; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_82; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_83; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_84; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_85; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_86; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_87; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_88; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_89; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_90; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_91; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_92; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_93; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_94; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_95; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_96; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_97; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_98; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_99; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_100; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_101; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_102; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_103; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_104; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_105; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_106; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_107; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_108; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_109; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_110; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_111; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_112; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_113; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_114; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_115; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_116; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_117; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_118; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_119; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_120; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_121; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_122; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_123; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_124; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_125; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_126; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_mask_127; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [8:0] u_rt_in_io_sc2mac_dat_pd; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_dat_pvld; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_1; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_2; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_3; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_4; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_5; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_6; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_7; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_8; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_9; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_10; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_11; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_12; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_13; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_14; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_15; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_16; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_17; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_18; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_19; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_20; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_21; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_22; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_23; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_24; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_25; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_26; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_27; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_28; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_29; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_30; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_31; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_32; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_33; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_34; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_35; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_36; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_37; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_38; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_39; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_40; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_41; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_42; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_43; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_44; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_45; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_46; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_47; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_48; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_49; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_50; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_51; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_52; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_53; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_54; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_55; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_56; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_57; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_58; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_59; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_60; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_61; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_62; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_63; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_64; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_65; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_66; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_67; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_68; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_69; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_70; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_71; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_72; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_73; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_74; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_75; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_76; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_77; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_78; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_79; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_80; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_81; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_82; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_83; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_84; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_85; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_86; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_87; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_88; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_89; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_90; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_91; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_92; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_93; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_94; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_95; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_96; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_97; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_98; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_99; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_100; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_101; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_102; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_103; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_104; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_105; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_106; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_107; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_108; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_109; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_110; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_111; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_112; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_113; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_114; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_115; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_116; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_117; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_118; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_119; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_120; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_121; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_122; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_123; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_124; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_125; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_126; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_sc2mac_wt_data_127; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_1; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_2; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_3; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_4; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_5; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_6; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_7; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_8; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_9; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_10; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_11; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_12; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_13; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_14; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_15; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_16; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_17; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_18; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_19; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_20; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_21; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_22; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_23; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_24; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_25; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_26; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_27; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_28; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_29; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_30; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_31; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_32; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_33; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_34; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_35; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_36; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_37; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_38; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_39; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_40; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_41; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_42; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_43; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_44; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_45; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_46; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_47; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_48; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_49; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_50; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_51; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_52; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_53; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_54; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_55; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_56; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_57; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_58; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_59; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_60; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_61; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_62; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_63; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_64; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_65; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_66; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_67; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_68; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_69; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_70; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_71; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_72; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_73; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_74; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_75; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_76; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_77; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_78; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_79; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_80; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_81; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_82; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_83; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_84; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_85; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_86; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_87; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_88; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_89; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_90; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_91; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_92; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_93; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_94; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_95; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_96; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_97; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_98; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_99; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_100; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_101; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_102; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_103; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_104; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_105; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_106; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_107; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_108; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_109; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_110; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_111; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_112; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_113; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_114; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_115; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_116; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_117; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_118; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_119; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_120; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_121; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_122; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_123; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_124; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_125; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_126; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_mask_127; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_sel_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_sc2mac_wt_pvld; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_1; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_2; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_3; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_4; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_5; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_6; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_7; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_8; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_9; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_10; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_11; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_12; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_13; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_14; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_15; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_16; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_17; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_18; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_19; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_20; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_21; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_22; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_23; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_24; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_25; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_26; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_27; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_28; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_29; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_30; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_31; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_32; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_33; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_34; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_35; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_36; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_37; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_38; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_39; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_40; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_41; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_42; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_43; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_44; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_45; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_46; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_47; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_48; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_49; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_50; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_51; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_52; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_53; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_54; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_55; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_56; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_57; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_58; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_59; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_60; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_61; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_62; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_63; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_64; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_65; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_66; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_67; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_68; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_69; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_70; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_71; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_72; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_73; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_74; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_75; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_76; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_77; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_78; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_79; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_80; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_81; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_82; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_83; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_84; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_85; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_86; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_87; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_88; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_89; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_90; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_91; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_92; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_93; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_94; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_95; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_96; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_97; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_98; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_99; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_100; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_101; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_102; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_103; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_104; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_105; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_106; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_107; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_108; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_109; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_110; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_111; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_112; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_113; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_114; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_115; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_116; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_117; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_118; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_119; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_120; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_121; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_122; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_123; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_124; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_125; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_126; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_dat_data_127; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_1; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_2; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_3; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_4; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_5; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_6; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_7; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_8; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_9; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_10; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_11; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_12; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_13; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_14; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_15; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_16; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_17; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_18; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_19; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_20; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_21; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_22; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_23; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_24; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_25; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_26; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_27; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_28; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_29; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_30; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_31; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_32; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_33; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_34; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_35; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_36; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_37; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_38; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_39; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_40; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_41; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_42; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_43; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_44; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_45; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_46; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_47; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_48; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_49; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_50; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_51; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_52; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_53; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_54; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_55; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_56; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_57; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_58; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_59; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_60; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_61; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_62; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_63; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_64; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_65; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_66; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_67; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_68; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_69; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_70; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_71; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_72; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_73; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_74; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_75; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_76; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_77; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_78; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_79; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_80; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_81; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_82; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_83; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_84; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_85; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_86; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_87; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_88; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_89; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_90; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_91; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_92; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_93; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_94; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_95; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_96; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_97; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_98; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_99; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_100; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_101; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_102; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_103; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_104; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_105; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_106; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_107; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_108; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_109; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_110; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_111; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_112; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_113; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_114; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_115; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_116; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_117; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_118; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_119; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_120; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_121; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_122; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_123; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_124; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_125; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_126; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_mask_127; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [8:0] u_rt_in_io_in_dat_pd; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_pvld; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_stripe_st; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_dat_stripe_end; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_1; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_2; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_3; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_4; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_5; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_6; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_7; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_8; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_9; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_10; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_11; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_12; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_13; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_14; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_15; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_16; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_17; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_18; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_19; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_20; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_21; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_22; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_23; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_24; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_25; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_26; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_27; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_28; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_29; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_30; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_31; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_32; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_33; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_34; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_35; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_36; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_37; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_38; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_39; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_40; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_41; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_42; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_43; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_44; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_45; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_46; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_47; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_48; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_49; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_50; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_51; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_52; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_53; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_54; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_55; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_56; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_57; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_58; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_59; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_60; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_61; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_62; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_63; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_64; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_65; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_66; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_67; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_68; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_69; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_70; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_71; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_72; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_73; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_74; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_75; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_76; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_77; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_78; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_79; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_80; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_81; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_82; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_83; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_84; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_85; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_86; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_87; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_88; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_89; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_90; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_91; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_92; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_93; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_94; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_95; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_96; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_97; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_98; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_99; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_100; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_101; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_102; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_103; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_104; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_105; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_106; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_107; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_108; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_109; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_110; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_111; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_112; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_113; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_114; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_115; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_116; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_117; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_118; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_119; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_120; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_121; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_122; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_123; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_124; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_125; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_126; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire [7:0] u_rt_in_io_in_wt_data_127; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_1; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_2; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_3; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_4; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_5; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_6; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_7; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_8; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_9; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_10; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_11; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_12; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_13; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_14; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_15; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_16; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_17; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_18; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_19; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_20; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_21; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_22; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_23; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_24; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_25; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_26; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_27; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_28; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_29; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_30; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_31; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_32; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_33; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_34; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_35; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_36; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_37; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_38; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_39; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_40; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_41; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_42; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_43; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_44; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_45; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_46; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_47; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_48; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_49; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_50; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_51; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_52; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_53; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_54; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_55; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_56; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_57; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_58; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_59; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_60; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_61; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_62; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_63; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_64; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_65; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_66; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_67; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_68; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_69; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_70; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_71; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_72; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_73; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_74; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_75; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_76; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_77; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_78; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_79; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_80; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_81; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_82; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_83; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_84; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_85; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_86; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_87; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_88; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_89; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_90; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_91; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_92; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_93; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_94; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_95; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_96; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_97; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_98; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_99; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_100; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_101; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_102; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_103; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_104; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_105; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_106; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_107; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_108; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_109; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_110; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_111; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_112; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_113; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_114; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_115; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_116; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_117; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_118; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_119; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_120; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_121; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_122; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_123; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_124; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_125; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_126; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_mask_127; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_sel_0; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_rt_in_io_in_wt_pvld; // @[NV_NVDLA_CMAC_core.scala 52:25]
  wire  u_active_clock; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_reset; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_dat_data_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_mask_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_pvld; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_stripe_st; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_dat_stripe_end; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_in_wt_data_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_mask_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_pvld; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_in_wt_sel_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_dat_actv_data_0_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_nz_0_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_dat_actv_pvld_0_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire [7:0] u_active_io_wt_actv_data_0_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_nz_0_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_0; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_1; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_2; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_3; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_4; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_5; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_6; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_7; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_8; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_9; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_10; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_11; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_12; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_13; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_14; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_15; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_16; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_17; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_18; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_19; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_20; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_21; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_22; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_23; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_24; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_25; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_26; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_27; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_28; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_29; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_30; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_31; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_32; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_33; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_34; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_35; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_36; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_37; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_38; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_39; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_40; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_41; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_42; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_43; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_44; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_45; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_46; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_47; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_48; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_49; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_50; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_51; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_52; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_53; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_54; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_55; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_56; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_57; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_58; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_59; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_60; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_61; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_62; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_63; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_64; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_65; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_66; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_67; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_68; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_69; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_70; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_71; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_72; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_73; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_74; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_75; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_76; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_77; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_78; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_79; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_80; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_81; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_82; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_83; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_84; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_85; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_86; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_87; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_88; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_89; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_90; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_91; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_92; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_93; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_94; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_95; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_96; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_97; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_98; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_99; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_100; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_101; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_102; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_103; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_104; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_105; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_106; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_107; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_108; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_109; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_110; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_111; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_112; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_113; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_114; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_115; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_116; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_117; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_118; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_119; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_120; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_121; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_122; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_123; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_124; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_125; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_126; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  u_active_io_wt_actv_pvld_0_127; // @[NV_NVDLA_CMAC_core.scala 82:26]
  wire  NV_NVDLA_CMAC_CORE_mac_clock; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_0; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_1; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_2; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_3; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_4; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_5; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_6; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_7; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_8; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_9; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_10; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_11; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_12; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_13; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_14; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_15; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_16; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_17; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_18; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_19; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_20; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_21; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_22; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_23; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_24; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_25; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_26; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_27; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_28; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_29; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_30; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_31; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_32; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_33; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_34; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_35; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_36; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_37; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_38; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_39; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_40; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_41; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_42; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_43; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_44; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_45; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_46; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_47; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_48; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_49; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_50; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_51; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_52; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_53; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_54; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_55; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_56; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_57; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_58; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_59; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_60; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_61; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_62; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_63; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_64; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_65; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_66; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_67; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_68; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_69; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_70; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_71; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_72; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_73; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_74; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_75; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_76; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_77; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_78; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_79; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_80; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_81; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_82; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_83; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_84; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_85; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_86; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_87; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_88; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_89; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_90; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_91; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_92; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_93; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_94; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_95; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_96; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_97; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_98; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_99; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_100; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_101; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_102; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_103; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_104; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_105; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_106; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_107; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_108; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_109; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_110; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_111; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_112; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_113; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_114; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_115; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_116; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_117; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_118; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_119; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_120; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_121; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_122; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_123; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_124; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_125; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_126; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_127; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_0; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_1; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_2; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_3; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_4; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_5; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_6; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_7; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_8; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_9; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_10; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_11; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_12; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_13; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_14; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_15; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_16; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_17; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_18; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_19; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_20; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_21; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_22; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_23; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_24; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_25; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_26; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_27; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_28; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_29; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_30; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_31; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_32; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_33; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_34; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_35; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_36; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_37; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_38; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_39; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_40; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_41; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_42; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_43; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_44; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_45; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_46; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_47; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_48; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_49; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_50; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_51; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_52; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_53; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_54; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_55; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_56; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_57; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_58; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_59; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_60; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_61; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_62; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_63; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_64; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_65; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_66; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_67; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_68; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_69; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_70; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_71; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_72; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_73; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_74; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_75; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_76; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_77; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_78; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_79; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_80; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_81; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_82; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_83; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_84; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_85; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_86; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_87; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_88; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_89; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_90; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_91; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_92; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_93; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_94; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_95; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_96; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_97; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_98; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_99; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_100; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_101; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_102; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_103; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_104; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_105; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_106; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_107; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_108; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_109; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_110; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_111; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_112; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_113; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_114; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_115; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_116; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_117; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_118; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_119; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_120; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_121; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_122; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_123; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_124; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_125; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_126; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_127; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_0; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_1; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_2; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_3; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_4; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_5; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_6; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_7; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_8; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_9; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_10; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_11; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_12; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_13; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_14; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_15; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_16; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_17; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_18; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_19; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_20; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_21; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_22; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_23; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_24; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_25; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_26; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_27; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_28; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_29; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_30; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_31; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_32; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_33; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_34; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_35; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_36; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_37; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_38; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_39; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_40; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_41; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_42; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_43; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_44; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_45; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_46; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_47; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_48; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_49; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_50; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_51; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_52; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_53; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_54; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_55; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_56; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_57; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_58; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_59; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_60; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_61; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_62; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_63; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_64; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_65; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_66; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_67; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_68; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_69; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_70; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_71; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_72; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_73; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_74; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_75; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_76; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_77; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_78; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_79; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_80; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_81; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_82; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_83; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_84; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_85; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_86; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_87; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_88; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_89; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_90; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_91; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_92; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_93; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_94; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_95; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_96; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_97; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_98; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_99; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_100; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_101; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_102; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_103; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_104; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_105; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_106; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_107; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_108; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_109; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_110; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_111; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_112; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_113; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_114; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_115; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_116; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_117; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_118; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_119; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_120; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_121; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_122; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_123; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_124; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_125; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_126; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_127; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_0; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_1; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_2; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_3; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_4; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_5; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_6; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_7; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_8; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_9; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_10; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_11; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_12; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_13; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_14; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_15; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_16; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_17; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_18; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_19; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_20; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_21; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_22; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_23; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_24; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_25; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_26; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_27; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_28; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_29; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_30; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_31; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_32; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_33; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_34; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_35; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_36; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_37; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_38; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_39; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_40; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_41; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_42; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_43; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_44; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_45; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_46; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_47; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_48; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_49; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_50; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_51; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_52; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_53; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_54; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_55; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_56; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_57; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_58; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_59; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_60; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_61; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_62; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_63; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_64; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_65; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_66; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_67; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_68; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_69; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_70; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_71; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_72; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_73; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_74; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_75; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_76; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_77; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_78; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_79; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_80; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_81; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_82; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_83; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_84; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_85; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_86; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_87; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_88; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_89; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_90; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_91; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_92; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_93; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_94; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_95; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_96; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_97; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_98; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_99; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_100; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_101; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_102; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_103; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_104; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_105; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_106; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_107; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_108; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_109; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_110; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_111; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_112; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_113; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_114; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_115; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_116; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_117; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_118; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_119; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_120; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_121; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_122; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_123; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_124; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_125; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_126; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [7:0] NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_127; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_0; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_1; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_2; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_3; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_4; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_5; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_6; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_7; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_8; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_9; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_10; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_11; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_12; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_13; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_14; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_15; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_16; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_17; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_18; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_19; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_20; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_21; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_22; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_23; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_24; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_25; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_26; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_27; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_28; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_29; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_30; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_31; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_32; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_33; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_34; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_35; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_36; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_37; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_38; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_39; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_40; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_41; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_42; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_43; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_44; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_45; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_46; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_47; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_48; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_49; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_50; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_51; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_52; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_53; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_54; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_55; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_56; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_57; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_58; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_59; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_60; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_61; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_62; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_63; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_64; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_65; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_66; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_67; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_68; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_69; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_70; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_71; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_72; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_73; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_74; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_75; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_76; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_77; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_78; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_79; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_80; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_81; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_82; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_83; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_84; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_85; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_86; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_87; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_88; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_89; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_90; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_91; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_92; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_93; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_94; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_95; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_96; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_97; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_98; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_99; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_100; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_101; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_102; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_103; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_104; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_105; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_106; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_107; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_108; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_109; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_110; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_111; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_112; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_113; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_114; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_115; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_116; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_117; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_118; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_119; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_120; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_121; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_122; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_123; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_124; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_125; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_126; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_127; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_0; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_1; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_2; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_3; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_4; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_5; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_6; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_7; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_8; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_9; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_10; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_11; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_12; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_13; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_14; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_15; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_16; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_17; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_18; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_19; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_20; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_21; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_22; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_23; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_24; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_25; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_26; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_27; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_28; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_29; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_30; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_31; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_32; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_33; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_34; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_35; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_36; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_37; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_38; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_39; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_40; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_41; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_42; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_43; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_44; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_45; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_46; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_47; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_48; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_49; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_50; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_51; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_52; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_53; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_54; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_55; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_56; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_57; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_58; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_59; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_60; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_61; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_62; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_63; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_64; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_65; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_66; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_67; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_68; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_69; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_70; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_71; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_72; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_73; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_74; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_75; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_76; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_77; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_78; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_79; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_80; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_81; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_82; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_83; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_84; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_85; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_86; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_87; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_88; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_89; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_90; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_91; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_92; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_93; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_94; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_95; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_96; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_97; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_98; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_99; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_100; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_101; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_102; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_103; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_104; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_105; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_106; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_107; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_108; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_109; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_110; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_111; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_112; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_113; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_114; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_115; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_116; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_117; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_118; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_119; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_120; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_121; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_122; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_123; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_124; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_125; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_126; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_127; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire [22:0] NV_NVDLA_CMAC_CORE_mac_io_mac_out_data; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  NV_NVDLA_CMAC_CORE_mac_io_mac_out_pvld; // @[NV_NVDLA_CMAC_core.scala 108:56]
  wire  u_rt_out_clock; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire  u_rt_out_reset; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire [22:0] u_rt_out_io_out_data_0; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire  u_rt_out_io_out_mask_0; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire [8:0] u_rt_out_io_out_pd; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire  u_rt_out_io_out_pvld; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire [22:0] u_rt_out_io_mac2accu_data_0; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire  u_rt_out_io_mac2accu_mask_0; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire [8:0] u_rt_out_io_mac2accu_pd; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire  u_rt_out_io_mac2accu_pvld; // @[NV_NVDLA_CMAC_core.scala 129:26]
  wire  u_rt_out_io_dp2reg_done; // @[NV_NVDLA_CMAC_core.scala 129:26]
  reg  _T_1119; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  reg  out_pvld; // @[Reg.scala 11:16]
  reg [31:0] _RAND_1;
  reg [8:0] _T_1122; // @[Reg.scala 11:16]
  reg [31:0] _RAND_2;
  reg [8:0] out_pd; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  NV_NVDLA_CMAC_CORE_rt_in u_rt_in ( // @[NV_NVDLA_CMAC_core.scala 52:25]
    .clock(u_rt_in_clock),
    .reset(u_rt_in_reset),
    .io_sc2mac_dat_data_0(u_rt_in_io_sc2mac_dat_data_0),
    .io_sc2mac_dat_data_1(u_rt_in_io_sc2mac_dat_data_1),
    .io_sc2mac_dat_data_2(u_rt_in_io_sc2mac_dat_data_2),
    .io_sc2mac_dat_data_3(u_rt_in_io_sc2mac_dat_data_3),
    .io_sc2mac_dat_data_4(u_rt_in_io_sc2mac_dat_data_4),
    .io_sc2mac_dat_data_5(u_rt_in_io_sc2mac_dat_data_5),
    .io_sc2mac_dat_data_6(u_rt_in_io_sc2mac_dat_data_6),
    .io_sc2mac_dat_data_7(u_rt_in_io_sc2mac_dat_data_7),
    .io_sc2mac_dat_data_8(u_rt_in_io_sc2mac_dat_data_8),
    .io_sc2mac_dat_data_9(u_rt_in_io_sc2mac_dat_data_9),
    .io_sc2mac_dat_data_10(u_rt_in_io_sc2mac_dat_data_10),
    .io_sc2mac_dat_data_11(u_rt_in_io_sc2mac_dat_data_11),
    .io_sc2mac_dat_data_12(u_rt_in_io_sc2mac_dat_data_12),
    .io_sc2mac_dat_data_13(u_rt_in_io_sc2mac_dat_data_13),
    .io_sc2mac_dat_data_14(u_rt_in_io_sc2mac_dat_data_14),
    .io_sc2mac_dat_data_15(u_rt_in_io_sc2mac_dat_data_15),
    .io_sc2mac_dat_data_16(u_rt_in_io_sc2mac_dat_data_16),
    .io_sc2mac_dat_data_17(u_rt_in_io_sc2mac_dat_data_17),
    .io_sc2mac_dat_data_18(u_rt_in_io_sc2mac_dat_data_18),
    .io_sc2mac_dat_data_19(u_rt_in_io_sc2mac_dat_data_19),
    .io_sc2mac_dat_data_20(u_rt_in_io_sc2mac_dat_data_20),
    .io_sc2mac_dat_data_21(u_rt_in_io_sc2mac_dat_data_21),
    .io_sc2mac_dat_data_22(u_rt_in_io_sc2mac_dat_data_22),
    .io_sc2mac_dat_data_23(u_rt_in_io_sc2mac_dat_data_23),
    .io_sc2mac_dat_data_24(u_rt_in_io_sc2mac_dat_data_24),
    .io_sc2mac_dat_data_25(u_rt_in_io_sc2mac_dat_data_25),
    .io_sc2mac_dat_data_26(u_rt_in_io_sc2mac_dat_data_26),
    .io_sc2mac_dat_data_27(u_rt_in_io_sc2mac_dat_data_27),
    .io_sc2mac_dat_data_28(u_rt_in_io_sc2mac_dat_data_28),
    .io_sc2mac_dat_data_29(u_rt_in_io_sc2mac_dat_data_29),
    .io_sc2mac_dat_data_30(u_rt_in_io_sc2mac_dat_data_30),
    .io_sc2mac_dat_data_31(u_rt_in_io_sc2mac_dat_data_31),
    .io_sc2mac_dat_data_32(u_rt_in_io_sc2mac_dat_data_32),
    .io_sc2mac_dat_data_33(u_rt_in_io_sc2mac_dat_data_33),
    .io_sc2mac_dat_data_34(u_rt_in_io_sc2mac_dat_data_34),
    .io_sc2mac_dat_data_35(u_rt_in_io_sc2mac_dat_data_35),
    .io_sc2mac_dat_data_36(u_rt_in_io_sc2mac_dat_data_36),
    .io_sc2mac_dat_data_37(u_rt_in_io_sc2mac_dat_data_37),
    .io_sc2mac_dat_data_38(u_rt_in_io_sc2mac_dat_data_38),
    .io_sc2mac_dat_data_39(u_rt_in_io_sc2mac_dat_data_39),
    .io_sc2mac_dat_data_40(u_rt_in_io_sc2mac_dat_data_40),
    .io_sc2mac_dat_data_41(u_rt_in_io_sc2mac_dat_data_41),
    .io_sc2mac_dat_data_42(u_rt_in_io_sc2mac_dat_data_42),
    .io_sc2mac_dat_data_43(u_rt_in_io_sc2mac_dat_data_43),
    .io_sc2mac_dat_data_44(u_rt_in_io_sc2mac_dat_data_44),
    .io_sc2mac_dat_data_45(u_rt_in_io_sc2mac_dat_data_45),
    .io_sc2mac_dat_data_46(u_rt_in_io_sc2mac_dat_data_46),
    .io_sc2mac_dat_data_47(u_rt_in_io_sc2mac_dat_data_47),
    .io_sc2mac_dat_data_48(u_rt_in_io_sc2mac_dat_data_48),
    .io_sc2mac_dat_data_49(u_rt_in_io_sc2mac_dat_data_49),
    .io_sc2mac_dat_data_50(u_rt_in_io_sc2mac_dat_data_50),
    .io_sc2mac_dat_data_51(u_rt_in_io_sc2mac_dat_data_51),
    .io_sc2mac_dat_data_52(u_rt_in_io_sc2mac_dat_data_52),
    .io_sc2mac_dat_data_53(u_rt_in_io_sc2mac_dat_data_53),
    .io_sc2mac_dat_data_54(u_rt_in_io_sc2mac_dat_data_54),
    .io_sc2mac_dat_data_55(u_rt_in_io_sc2mac_dat_data_55),
    .io_sc2mac_dat_data_56(u_rt_in_io_sc2mac_dat_data_56),
    .io_sc2mac_dat_data_57(u_rt_in_io_sc2mac_dat_data_57),
    .io_sc2mac_dat_data_58(u_rt_in_io_sc2mac_dat_data_58),
    .io_sc2mac_dat_data_59(u_rt_in_io_sc2mac_dat_data_59),
    .io_sc2mac_dat_data_60(u_rt_in_io_sc2mac_dat_data_60),
    .io_sc2mac_dat_data_61(u_rt_in_io_sc2mac_dat_data_61),
    .io_sc2mac_dat_data_62(u_rt_in_io_sc2mac_dat_data_62),
    .io_sc2mac_dat_data_63(u_rt_in_io_sc2mac_dat_data_63),
    .io_sc2mac_dat_data_64(u_rt_in_io_sc2mac_dat_data_64),
    .io_sc2mac_dat_data_65(u_rt_in_io_sc2mac_dat_data_65),
    .io_sc2mac_dat_data_66(u_rt_in_io_sc2mac_dat_data_66),
    .io_sc2mac_dat_data_67(u_rt_in_io_sc2mac_dat_data_67),
    .io_sc2mac_dat_data_68(u_rt_in_io_sc2mac_dat_data_68),
    .io_sc2mac_dat_data_69(u_rt_in_io_sc2mac_dat_data_69),
    .io_sc2mac_dat_data_70(u_rt_in_io_sc2mac_dat_data_70),
    .io_sc2mac_dat_data_71(u_rt_in_io_sc2mac_dat_data_71),
    .io_sc2mac_dat_data_72(u_rt_in_io_sc2mac_dat_data_72),
    .io_sc2mac_dat_data_73(u_rt_in_io_sc2mac_dat_data_73),
    .io_sc2mac_dat_data_74(u_rt_in_io_sc2mac_dat_data_74),
    .io_sc2mac_dat_data_75(u_rt_in_io_sc2mac_dat_data_75),
    .io_sc2mac_dat_data_76(u_rt_in_io_sc2mac_dat_data_76),
    .io_sc2mac_dat_data_77(u_rt_in_io_sc2mac_dat_data_77),
    .io_sc2mac_dat_data_78(u_rt_in_io_sc2mac_dat_data_78),
    .io_sc2mac_dat_data_79(u_rt_in_io_sc2mac_dat_data_79),
    .io_sc2mac_dat_data_80(u_rt_in_io_sc2mac_dat_data_80),
    .io_sc2mac_dat_data_81(u_rt_in_io_sc2mac_dat_data_81),
    .io_sc2mac_dat_data_82(u_rt_in_io_sc2mac_dat_data_82),
    .io_sc2mac_dat_data_83(u_rt_in_io_sc2mac_dat_data_83),
    .io_sc2mac_dat_data_84(u_rt_in_io_sc2mac_dat_data_84),
    .io_sc2mac_dat_data_85(u_rt_in_io_sc2mac_dat_data_85),
    .io_sc2mac_dat_data_86(u_rt_in_io_sc2mac_dat_data_86),
    .io_sc2mac_dat_data_87(u_rt_in_io_sc2mac_dat_data_87),
    .io_sc2mac_dat_data_88(u_rt_in_io_sc2mac_dat_data_88),
    .io_sc2mac_dat_data_89(u_rt_in_io_sc2mac_dat_data_89),
    .io_sc2mac_dat_data_90(u_rt_in_io_sc2mac_dat_data_90),
    .io_sc2mac_dat_data_91(u_rt_in_io_sc2mac_dat_data_91),
    .io_sc2mac_dat_data_92(u_rt_in_io_sc2mac_dat_data_92),
    .io_sc2mac_dat_data_93(u_rt_in_io_sc2mac_dat_data_93),
    .io_sc2mac_dat_data_94(u_rt_in_io_sc2mac_dat_data_94),
    .io_sc2mac_dat_data_95(u_rt_in_io_sc2mac_dat_data_95),
    .io_sc2mac_dat_data_96(u_rt_in_io_sc2mac_dat_data_96),
    .io_sc2mac_dat_data_97(u_rt_in_io_sc2mac_dat_data_97),
    .io_sc2mac_dat_data_98(u_rt_in_io_sc2mac_dat_data_98),
    .io_sc2mac_dat_data_99(u_rt_in_io_sc2mac_dat_data_99),
    .io_sc2mac_dat_data_100(u_rt_in_io_sc2mac_dat_data_100),
    .io_sc2mac_dat_data_101(u_rt_in_io_sc2mac_dat_data_101),
    .io_sc2mac_dat_data_102(u_rt_in_io_sc2mac_dat_data_102),
    .io_sc2mac_dat_data_103(u_rt_in_io_sc2mac_dat_data_103),
    .io_sc2mac_dat_data_104(u_rt_in_io_sc2mac_dat_data_104),
    .io_sc2mac_dat_data_105(u_rt_in_io_sc2mac_dat_data_105),
    .io_sc2mac_dat_data_106(u_rt_in_io_sc2mac_dat_data_106),
    .io_sc2mac_dat_data_107(u_rt_in_io_sc2mac_dat_data_107),
    .io_sc2mac_dat_data_108(u_rt_in_io_sc2mac_dat_data_108),
    .io_sc2mac_dat_data_109(u_rt_in_io_sc2mac_dat_data_109),
    .io_sc2mac_dat_data_110(u_rt_in_io_sc2mac_dat_data_110),
    .io_sc2mac_dat_data_111(u_rt_in_io_sc2mac_dat_data_111),
    .io_sc2mac_dat_data_112(u_rt_in_io_sc2mac_dat_data_112),
    .io_sc2mac_dat_data_113(u_rt_in_io_sc2mac_dat_data_113),
    .io_sc2mac_dat_data_114(u_rt_in_io_sc2mac_dat_data_114),
    .io_sc2mac_dat_data_115(u_rt_in_io_sc2mac_dat_data_115),
    .io_sc2mac_dat_data_116(u_rt_in_io_sc2mac_dat_data_116),
    .io_sc2mac_dat_data_117(u_rt_in_io_sc2mac_dat_data_117),
    .io_sc2mac_dat_data_118(u_rt_in_io_sc2mac_dat_data_118),
    .io_sc2mac_dat_data_119(u_rt_in_io_sc2mac_dat_data_119),
    .io_sc2mac_dat_data_120(u_rt_in_io_sc2mac_dat_data_120),
    .io_sc2mac_dat_data_121(u_rt_in_io_sc2mac_dat_data_121),
    .io_sc2mac_dat_data_122(u_rt_in_io_sc2mac_dat_data_122),
    .io_sc2mac_dat_data_123(u_rt_in_io_sc2mac_dat_data_123),
    .io_sc2mac_dat_data_124(u_rt_in_io_sc2mac_dat_data_124),
    .io_sc2mac_dat_data_125(u_rt_in_io_sc2mac_dat_data_125),
    .io_sc2mac_dat_data_126(u_rt_in_io_sc2mac_dat_data_126),
    .io_sc2mac_dat_data_127(u_rt_in_io_sc2mac_dat_data_127),
    .io_sc2mac_dat_mask_0(u_rt_in_io_sc2mac_dat_mask_0),
    .io_sc2mac_dat_mask_1(u_rt_in_io_sc2mac_dat_mask_1),
    .io_sc2mac_dat_mask_2(u_rt_in_io_sc2mac_dat_mask_2),
    .io_sc2mac_dat_mask_3(u_rt_in_io_sc2mac_dat_mask_3),
    .io_sc2mac_dat_mask_4(u_rt_in_io_sc2mac_dat_mask_4),
    .io_sc2mac_dat_mask_5(u_rt_in_io_sc2mac_dat_mask_5),
    .io_sc2mac_dat_mask_6(u_rt_in_io_sc2mac_dat_mask_6),
    .io_sc2mac_dat_mask_7(u_rt_in_io_sc2mac_dat_mask_7),
    .io_sc2mac_dat_mask_8(u_rt_in_io_sc2mac_dat_mask_8),
    .io_sc2mac_dat_mask_9(u_rt_in_io_sc2mac_dat_mask_9),
    .io_sc2mac_dat_mask_10(u_rt_in_io_sc2mac_dat_mask_10),
    .io_sc2mac_dat_mask_11(u_rt_in_io_sc2mac_dat_mask_11),
    .io_sc2mac_dat_mask_12(u_rt_in_io_sc2mac_dat_mask_12),
    .io_sc2mac_dat_mask_13(u_rt_in_io_sc2mac_dat_mask_13),
    .io_sc2mac_dat_mask_14(u_rt_in_io_sc2mac_dat_mask_14),
    .io_sc2mac_dat_mask_15(u_rt_in_io_sc2mac_dat_mask_15),
    .io_sc2mac_dat_mask_16(u_rt_in_io_sc2mac_dat_mask_16),
    .io_sc2mac_dat_mask_17(u_rt_in_io_sc2mac_dat_mask_17),
    .io_sc2mac_dat_mask_18(u_rt_in_io_sc2mac_dat_mask_18),
    .io_sc2mac_dat_mask_19(u_rt_in_io_sc2mac_dat_mask_19),
    .io_sc2mac_dat_mask_20(u_rt_in_io_sc2mac_dat_mask_20),
    .io_sc2mac_dat_mask_21(u_rt_in_io_sc2mac_dat_mask_21),
    .io_sc2mac_dat_mask_22(u_rt_in_io_sc2mac_dat_mask_22),
    .io_sc2mac_dat_mask_23(u_rt_in_io_sc2mac_dat_mask_23),
    .io_sc2mac_dat_mask_24(u_rt_in_io_sc2mac_dat_mask_24),
    .io_sc2mac_dat_mask_25(u_rt_in_io_sc2mac_dat_mask_25),
    .io_sc2mac_dat_mask_26(u_rt_in_io_sc2mac_dat_mask_26),
    .io_sc2mac_dat_mask_27(u_rt_in_io_sc2mac_dat_mask_27),
    .io_sc2mac_dat_mask_28(u_rt_in_io_sc2mac_dat_mask_28),
    .io_sc2mac_dat_mask_29(u_rt_in_io_sc2mac_dat_mask_29),
    .io_sc2mac_dat_mask_30(u_rt_in_io_sc2mac_dat_mask_30),
    .io_sc2mac_dat_mask_31(u_rt_in_io_sc2mac_dat_mask_31),
    .io_sc2mac_dat_mask_32(u_rt_in_io_sc2mac_dat_mask_32),
    .io_sc2mac_dat_mask_33(u_rt_in_io_sc2mac_dat_mask_33),
    .io_sc2mac_dat_mask_34(u_rt_in_io_sc2mac_dat_mask_34),
    .io_sc2mac_dat_mask_35(u_rt_in_io_sc2mac_dat_mask_35),
    .io_sc2mac_dat_mask_36(u_rt_in_io_sc2mac_dat_mask_36),
    .io_sc2mac_dat_mask_37(u_rt_in_io_sc2mac_dat_mask_37),
    .io_sc2mac_dat_mask_38(u_rt_in_io_sc2mac_dat_mask_38),
    .io_sc2mac_dat_mask_39(u_rt_in_io_sc2mac_dat_mask_39),
    .io_sc2mac_dat_mask_40(u_rt_in_io_sc2mac_dat_mask_40),
    .io_sc2mac_dat_mask_41(u_rt_in_io_sc2mac_dat_mask_41),
    .io_sc2mac_dat_mask_42(u_rt_in_io_sc2mac_dat_mask_42),
    .io_sc2mac_dat_mask_43(u_rt_in_io_sc2mac_dat_mask_43),
    .io_sc2mac_dat_mask_44(u_rt_in_io_sc2mac_dat_mask_44),
    .io_sc2mac_dat_mask_45(u_rt_in_io_sc2mac_dat_mask_45),
    .io_sc2mac_dat_mask_46(u_rt_in_io_sc2mac_dat_mask_46),
    .io_sc2mac_dat_mask_47(u_rt_in_io_sc2mac_dat_mask_47),
    .io_sc2mac_dat_mask_48(u_rt_in_io_sc2mac_dat_mask_48),
    .io_sc2mac_dat_mask_49(u_rt_in_io_sc2mac_dat_mask_49),
    .io_sc2mac_dat_mask_50(u_rt_in_io_sc2mac_dat_mask_50),
    .io_sc2mac_dat_mask_51(u_rt_in_io_sc2mac_dat_mask_51),
    .io_sc2mac_dat_mask_52(u_rt_in_io_sc2mac_dat_mask_52),
    .io_sc2mac_dat_mask_53(u_rt_in_io_sc2mac_dat_mask_53),
    .io_sc2mac_dat_mask_54(u_rt_in_io_sc2mac_dat_mask_54),
    .io_sc2mac_dat_mask_55(u_rt_in_io_sc2mac_dat_mask_55),
    .io_sc2mac_dat_mask_56(u_rt_in_io_sc2mac_dat_mask_56),
    .io_sc2mac_dat_mask_57(u_rt_in_io_sc2mac_dat_mask_57),
    .io_sc2mac_dat_mask_58(u_rt_in_io_sc2mac_dat_mask_58),
    .io_sc2mac_dat_mask_59(u_rt_in_io_sc2mac_dat_mask_59),
    .io_sc2mac_dat_mask_60(u_rt_in_io_sc2mac_dat_mask_60),
    .io_sc2mac_dat_mask_61(u_rt_in_io_sc2mac_dat_mask_61),
    .io_sc2mac_dat_mask_62(u_rt_in_io_sc2mac_dat_mask_62),
    .io_sc2mac_dat_mask_63(u_rt_in_io_sc2mac_dat_mask_63),
    .io_sc2mac_dat_mask_64(u_rt_in_io_sc2mac_dat_mask_64),
    .io_sc2mac_dat_mask_65(u_rt_in_io_sc2mac_dat_mask_65),
    .io_sc2mac_dat_mask_66(u_rt_in_io_sc2mac_dat_mask_66),
    .io_sc2mac_dat_mask_67(u_rt_in_io_sc2mac_dat_mask_67),
    .io_sc2mac_dat_mask_68(u_rt_in_io_sc2mac_dat_mask_68),
    .io_sc2mac_dat_mask_69(u_rt_in_io_sc2mac_dat_mask_69),
    .io_sc2mac_dat_mask_70(u_rt_in_io_sc2mac_dat_mask_70),
    .io_sc2mac_dat_mask_71(u_rt_in_io_sc2mac_dat_mask_71),
    .io_sc2mac_dat_mask_72(u_rt_in_io_sc2mac_dat_mask_72),
    .io_sc2mac_dat_mask_73(u_rt_in_io_sc2mac_dat_mask_73),
    .io_sc2mac_dat_mask_74(u_rt_in_io_sc2mac_dat_mask_74),
    .io_sc2mac_dat_mask_75(u_rt_in_io_sc2mac_dat_mask_75),
    .io_sc2mac_dat_mask_76(u_rt_in_io_sc2mac_dat_mask_76),
    .io_sc2mac_dat_mask_77(u_rt_in_io_sc2mac_dat_mask_77),
    .io_sc2mac_dat_mask_78(u_rt_in_io_sc2mac_dat_mask_78),
    .io_sc2mac_dat_mask_79(u_rt_in_io_sc2mac_dat_mask_79),
    .io_sc2mac_dat_mask_80(u_rt_in_io_sc2mac_dat_mask_80),
    .io_sc2mac_dat_mask_81(u_rt_in_io_sc2mac_dat_mask_81),
    .io_sc2mac_dat_mask_82(u_rt_in_io_sc2mac_dat_mask_82),
    .io_sc2mac_dat_mask_83(u_rt_in_io_sc2mac_dat_mask_83),
    .io_sc2mac_dat_mask_84(u_rt_in_io_sc2mac_dat_mask_84),
    .io_sc2mac_dat_mask_85(u_rt_in_io_sc2mac_dat_mask_85),
    .io_sc2mac_dat_mask_86(u_rt_in_io_sc2mac_dat_mask_86),
    .io_sc2mac_dat_mask_87(u_rt_in_io_sc2mac_dat_mask_87),
    .io_sc2mac_dat_mask_88(u_rt_in_io_sc2mac_dat_mask_88),
    .io_sc2mac_dat_mask_89(u_rt_in_io_sc2mac_dat_mask_89),
    .io_sc2mac_dat_mask_90(u_rt_in_io_sc2mac_dat_mask_90),
    .io_sc2mac_dat_mask_91(u_rt_in_io_sc2mac_dat_mask_91),
    .io_sc2mac_dat_mask_92(u_rt_in_io_sc2mac_dat_mask_92),
    .io_sc2mac_dat_mask_93(u_rt_in_io_sc2mac_dat_mask_93),
    .io_sc2mac_dat_mask_94(u_rt_in_io_sc2mac_dat_mask_94),
    .io_sc2mac_dat_mask_95(u_rt_in_io_sc2mac_dat_mask_95),
    .io_sc2mac_dat_mask_96(u_rt_in_io_sc2mac_dat_mask_96),
    .io_sc2mac_dat_mask_97(u_rt_in_io_sc2mac_dat_mask_97),
    .io_sc2mac_dat_mask_98(u_rt_in_io_sc2mac_dat_mask_98),
    .io_sc2mac_dat_mask_99(u_rt_in_io_sc2mac_dat_mask_99),
    .io_sc2mac_dat_mask_100(u_rt_in_io_sc2mac_dat_mask_100),
    .io_sc2mac_dat_mask_101(u_rt_in_io_sc2mac_dat_mask_101),
    .io_sc2mac_dat_mask_102(u_rt_in_io_sc2mac_dat_mask_102),
    .io_sc2mac_dat_mask_103(u_rt_in_io_sc2mac_dat_mask_103),
    .io_sc2mac_dat_mask_104(u_rt_in_io_sc2mac_dat_mask_104),
    .io_sc2mac_dat_mask_105(u_rt_in_io_sc2mac_dat_mask_105),
    .io_sc2mac_dat_mask_106(u_rt_in_io_sc2mac_dat_mask_106),
    .io_sc2mac_dat_mask_107(u_rt_in_io_sc2mac_dat_mask_107),
    .io_sc2mac_dat_mask_108(u_rt_in_io_sc2mac_dat_mask_108),
    .io_sc2mac_dat_mask_109(u_rt_in_io_sc2mac_dat_mask_109),
    .io_sc2mac_dat_mask_110(u_rt_in_io_sc2mac_dat_mask_110),
    .io_sc2mac_dat_mask_111(u_rt_in_io_sc2mac_dat_mask_111),
    .io_sc2mac_dat_mask_112(u_rt_in_io_sc2mac_dat_mask_112),
    .io_sc2mac_dat_mask_113(u_rt_in_io_sc2mac_dat_mask_113),
    .io_sc2mac_dat_mask_114(u_rt_in_io_sc2mac_dat_mask_114),
    .io_sc2mac_dat_mask_115(u_rt_in_io_sc2mac_dat_mask_115),
    .io_sc2mac_dat_mask_116(u_rt_in_io_sc2mac_dat_mask_116),
    .io_sc2mac_dat_mask_117(u_rt_in_io_sc2mac_dat_mask_117),
    .io_sc2mac_dat_mask_118(u_rt_in_io_sc2mac_dat_mask_118),
    .io_sc2mac_dat_mask_119(u_rt_in_io_sc2mac_dat_mask_119),
    .io_sc2mac_dat_mask_120(u_rt_in_io_sc2mac_dat_mask_120),
    .io_sc2mac_dat_mask_121(u_rt_in_io_sc2mac_dat_mask_121),
    .io_sc2mac_dat_mask_122(u_rt_in_io_sc2mac_dat_mask_122),
    .io_sc2mac_dat_mask_123(u_rt_in_io_sc2mac_dat_mask_123),
    .io_sc2mac_dat_mask_124(u_rt_in_io_sc2mac_dat_mask_124),
    .io_sc2mac_dat_mask_125(u_rt_in_io_sc2mac_dat_mask_125),
    .io_sc2mac_dat_mask_126(u_rt_in_io_sc2mac_dat_mask_126),
    .io_sc2mac_dat_mask_127(u_rt_in_io_sc2mac_dat_mask_127),
    .io_sc2mac_dat_pd(u_rt_in_io_sc2mac_dat_pd),
    .io_sc2mac_dat_pvld(u_rt_in_io_sc2mac_dat_pvld),
    .io_sc2mac_wt_data_0(u_rt_in_io_sc2mac_wt_data_0),
    .io_sc2mac_wt_data_1(u_rt_in_io_sc2mac_wt_data_1),
    .io_sc2mac_wt_data_2(u_rt_in_io_sc2mac_wt_data_2),
    .io_sc2mac_wt_data_3(u_rt_in_io_sc2mac_wt_data_3),
    .io_sc2mac_wt_data_4(u_rt_in_io_sc2mac_wt_data_4),
    .io_sc2mac_wt_data_5(u_rt_in_io_sc2mac_wt_data_5),
    .io_sc2mac_wt_data_6(u_rt_in_io_sc2mac_wt_data_6),
    .io_sc2mac_wt_data_7(u_rt_in_io_sc2mac_wt_data_7),
    .io_sc2mac_wt_data_8(u_rt_in_io_sc2mac_wt_data_8),
    .io_sc2mac_wt_data_9(u_rt_in_io_sc2mac_wt_data_9),
    .io_sc2mac_wt_data_10(u_rt_in_io_sc2mac_wt_data_10),
    .io_sc2mac_wt_data_11(u_rt_in_io_sc2mac_wt_data_11),
    .io_sc2mac_wt_data_12(u_rt_in_io_sc2mac_wt_data_12),
    .io_sc2mac_wt_data_13(u_rt_in_io_sc2mac_wt_data_13),
    .io_sc2mac_wt_data_14(u_rt_in_io_sc2mac_wt_data_14),
    .io_sc2mac_wt_data_15(u_rt_in_io_sc2mac_wt_data_15),
    .io_sc2mac_wt_data_16(u_rt_in_io_sc2mac_wt_data_16),
    .io_sc2mac_wt_data_17(u_rt_in_io_sc2mac_wt_data_17),
    .io_sc2mac_wt_data_18(u_rt_in_io_sc2mac_wt_data_18),
    .io_sc2mac_wt_data_19(u_rt_in_io_sc2mac_wt_data_19),
    .io_sc2mac_wt_data_20(u_rt_in_io_sc2mac_wt_data_20),
    .io_sc2mac_wt_data_21(u_rt_in_io_sc2mac_wt_data_21),
    .io_sc2mac_wt_data_22(u_rt_in_io_sc2mac_wt_data_22),
    .io_sc2mac_wt_data_23(u_rt_in_io_sc2mac_wt_data_23),
    .io_sc2mac_wt_data_24(u_rt_in_io_sc2mac_wt_data_24),
    .io_sc2mac_wt_data_25(u_rt_in_io_sc2mac_wt_data_25),
    .io_sc2mac_wt_data_26(u_rt_in_io_sc2mac_wt_data_26),
    .io_sc2mac_wt_data_27(u_rt_in_io_sc2mac_wt_data_27),
    .io_sc2mac_wt_data_28(u_rt_in_io_sc2mac_wt_data_28),
    .io_sc2mac_wt_data_29(u_rt_in_io_sc2mac_wt_data_29),
    .io_sc2mac_wt_data_30(u_rt_in_io_sc2mac_wt_data_30),
    .io_sc2mac_wt_data_31(u_rt_in_io_sc2mac_wt_data_31),
    .io_sc2mac_wt_data_32(u_rt_in_io_sc2mac_wt_data_32),
    .io_sc2mac_wt_data_33(u_rt_in_io_sc2mac_wt_data_33),
    .io_sc2mac_wt_data_34(u_rt_in_io_sc2mac_wt_data_34),
    .io_sc2mac_wt_data_35(u_rt_in_io_sc2mac_wt_data_35),
    .io_sc2mac_wt_data_36(u_rt_in_io_sc2mac_wt_data_36),
    .io_sc2mac_wt_data_37(u_rt_in_io_sc2mac_wt_data_37),
    .io_sc2mac_wt_data_38(u_rt_in_io_sc2mac_wt_data_38),
    .io_sc2mac_wt_data_39(u_rt_in_io_sc2mac_wt_data_39),
    .io_sc2mac_wt_data_40(u_rt_in_io_sc2mac_wt_data_40),
    .io_sc2mac_wt_data_41(u_rt_in_io_sc2mac_wt_data_41),
    .io_sc2mac_wt_data_42(u_rt_in_io_sc2mac_wt_data_42),
    .io_sc2mac_wt_data_43(u_rt_in_io_sc2mac_wt_data_43),
    .io_sc2mac_wt_data_44(u_rt_in_io_sc2mac_wt_data_44),
    .io_sc2mac_wt_data_45(u_rt_in_io_sc2mac_wt_data_45),
    .io_sc2mac_wt_data_46(u_rt_in_io_sc2mac_wt_data_46),
    .io_sc2mac_wt_data_47(u_rt_in_io_sc2mac_wt_data_47),
    .io_sc2mac_wt_data_48(u_rt_in_io_sc2mac_wt_data_48),
    .io_sc2mac_wt_data_49(u_rt_in_io_sc2mac_wt_data_49),
    .io_sc2mac_wt_data_50(u_rt_in_io_sc2mac_wt_data_50),
    .io_sc2mac_wt_data_51(u_rt_in_io_sc2mac_wt_data_51),
    .io_sc2mac_wt_data_52(u_rt_in_io_sc2mac_wt_data_52),
    .io_sc2mac_wt_data_53(u_rt_in_io_sc2mac_wt_data_53),
    .io_sc2mac_wt_data_54(u_rt_in_io_sc2mac_wt_data_54),
    .io_sc2mac_wt_data_55(u_rt_in_io_sc2mac_wt_data_55),
    .io_sc2mac_wt_data_56(u_rt_in_io_sc2mac_wt_data_56),
    .io_sc2mac_wt_data_57(u_rt_in_io_sc2mac_wt_data_57),
    .io_sc2mac_wt_data_58(u_rt_in_io_sc2mac_wt_data_58),
    .io_sc2mac_wt_data_59(u_rt_in_io_sc2mac_wt_data_59),
    .io_sc2mac_wt_data_60(u_rt_in_io_sc2mac_wt_data_60),
    .io_sc2mac_wt_data_61(u_rt_in_io_sc2mac_wt_data_61),
    .io_sc2mac_wt_data_62(u_rt_in_io_sc2mac_wt_data_62),
    .io_sc2mac_wt_data_63(u_rt_in_io_sc2mac_wt_data_63),
    .io_sc2mac_wt_data_64(u_rt_in_io_sc2mac_wt_data_64),
    .io_sc2mac_wt_data_65(u_rt_in_io_sc2mac_wt_data_65),
    .io_sc2mac_wt_data_66(u_rt_in_io_sc2mac_wt_data_66),
    .io_sc2mac_wt_data_67(u_rt_in_io_sc2mac_wt_data_67),
    .io_sc2mac_wt_data_68(u_rt_in_io_sc2mac_wt_data_68),
    .io_sc2mac_wt_data_69(u_rt_in_io_sc2mac_wt_data_69),
    .io_sc2mac_wt_data_70(u_rt_in_io_sc2mac_wt_data_70),
    .io_sc2mac_wt_data_71(u_rt_in_io_sc2mac_wt_data_71),
    .io_sc2mac_wt_data_72(u_rt_in_io_sc2mac_wt_data_72),
    .io_sc2mac_wt_data_73(u_rt_in_io_sc2mac_wt_data_73),
    .io_sc2mac_wt_data_74(u_rt_in_io_sc2mac_wt_data_74),
    .io_sc2mac_wt_data_75(u_rt_in_io_sc2mac_wt_data_75),
    .io_sc2mac_wt_data_76(u_rt_in_io_sc2mac_wt_data_76),
    .io_sc2mac_wt_data_77(u_rt_in_io_sc2mac_wt_data_77),
    .io_sc2mac_wt_data_78(u_rt_in_io_sc2mac_wt_data_78),
    .io_sc2mac_wt_data_79(u_rt_in_io_sc2mac_wt_data_79),
    .io_sc2mac_wt_data_80(u_rt_in_io_sc2mac_wt_data_80),
    .io_sc2mac_wt_data_81(u_rt_in_io_sc2mac_wt_data_81),
    .io_sc2mac_wt_data_82(u_rt_in_io_sc2mac_wt_data_82),
    .io_sc2mac_wt_data_83(u_rt_in_io_sc2mac_wt_data_83),
    .io_sc2mac_wt_data_84(u_rt_in_io_sc2mac_wt_data_84),
    .io_sc2mac_wt_data_85(u_rt_in_io_sc2mac_wt_data_85),
    .io_sc2mac_wt_data_86(u_rt_in_io_sc2mac_wt_data_86),
    .io_sc2mac_wt_data_87(u_rt_in_io_sc2mac_wt_data_87),
    .io_sc2mac_wt_data_88(u_rt_in_io_sc2mac_wt_data_88),
    .io_sc2mac_wt_data_89(u_rt_in_io_sc2mac_wt_data_89),
    .io_sc2mac_wt_data_90(u_rt_in_io_sc2mac_wt_data_90),
    .io_sc2mac_wt_data_91(u_rt_in_io_sc2mac_wt_data_91),
    .io_sc2mac_wt_data_92(u_rt_in_io_sc2mac_wt_data_92),
    .io_sc2mac_wt_data_93(u_rt_in_io_sc2mac_wt_data_93),
    .io_sc2mac_wt_data_94(u_rt_in_io_sc2mac_wt_data_94),
    .io_sc2mac_wt_data_95(u_rt_in_io_sc2mac_wt_data_95),
    .io_sc2mac_wt_data_96(u_rt_in_io_sc2mac_wt_data_96),
    .io_sc2mac_wt_data_97(u_rt_in_io_sc2mac_wt_data_97),
    .io_sc2mac_wt_data_98(u_rt_in_io_sc2mac_wt_data_98),
    .io_sc2mac_wt_data_99(u_rt_in_io_sc2mac_wt_data_99),
    .io_sc2mac_wt_data_100(u_rt_in_io_sc2mac_wt_data_100),
    .io_sc2mac_wt_data_101(u_rt_in_io_sc2mac_wt_data_101),
    .io_sc2mac_wt_data_102(u_rt_in_io_sc2mac_wt_data_102),
    .io_sc2mac_wt_data_103(u_rt_in_io_sc2mac_wt_data_103),
    .io_sc2mac_wt_data_104(u_rt_in_io_sc2mac_wt_data_104),
    .io_sc2mac_wt_data_105(u_rt_in_io_sc2mac_wt_data_105),
    .io_sc2mac_wt_data_106(u_rt_in_io_sc2mac_wt_data_106),
    .io_sc2mac_wt_data_107(u_rt_in_io_sc2mac_wt_data_107),
    .io_sc2mac_wt_data_108(u_rt_in_io_sc2mac_wt_data_108),
    .io_sc2mac_wt_data_109(u_rt_in_io_sc2mac_wt_data_109),
    .io_sc2mac_wt_data_110(u_rt_in_io_sc2mac_wt_data_110),
    .io_sc2mac_wt_data_111(u_rt_in_io_sc2mac_wt_data_111),
    .io_sc2mac_wt_data_112(u_rt_in_io_sc2mac_wt_data_112),
    .io_sc2mac_wt_data_113(u_rt_in_io_sc2mac_wt_data_113),
    .io_sc2mac_wt_data_114(u_rt_in_io_sc2mac_wt_data_114),
    .io_sc2mac_wt_data_115(u_rt_in_io_sc2mac_wt_data_115),
    .io_sc2mac_wt_data_116(u_rt_in_io_sc2mac_wt_data_116),
    .io_sc2mac_wt_data_117(u_rt_in_io_sc2mac_wt_data_117),
    .io_sc2mac_wt_data_118(u_rt_in_io_sc2mac_wt_data_118),
    .io_sc2mac_wt_data_119(u_rt_in_io_sc2mac_wt_data_119),
    .io_sc2mac_wt_data_120(u_rt_in_io_sc2mac_wt_data_120),
    .io_sc2mac_wt_data_121(u_rt_in_io_sc2mac_wt_data_121),
    .io_sc2mac_wt_data_122(u_rt_in_io_sc2mac_wt_data_122),
    .io_sc2mac_wt_data_123(u_rt_in_io_sc2mac_wt_data_123),
    .io_sc2mac_wt_data_124(u_rt_in_io_sc2mac_wt_data_124),
    .io_sc2mac_wt_data_125(u_rt_in_io_sc2mac_wt_data_125),
    .io_sc2mac_wt_data_126(u_rt_in_io_sc2mac_wt_data_126),
    .io_sc2mac_wt_data_127(u_rt_in_io_sc2mac_wt_data_127),
    .io_sc2mac_wt_mask_0(u_rt_in_io_sc2mac_wt_mask_0),
    .io_sc2mac_wt_mask_1(u_rt_in_io_sc2mac_wt_mask_1),
    .io_sc2mac_wt_mask_2(u_rt_in_io_sc2mac_wt_mask_2),
    .io_sc2mac_wt_mask_3(u_rt_in_io_sc2mac_wt_mask_3),
    .io_sc2mac_wt_mask_4(u_rt_in_io_sc2mac_wt_mask_4),
    .io_sc2mac_wt_mask_5(u_rt_in_io_sc2mac_wt_mask_5),
    .io_sc2mac_wt_mask_6(u_rt_in_io_sc2mac_wt_mask_6),
    .io_sc2mac_wt_mask_7(u_rt_in_io_sc2mac_wt_mask_7),
    .io_sc2mac_wt_mask_8(u_rt_in_io_sc2mac_wt_mask_8),
    .io_sc2mac_wt_mask_9(u_rt_in_io_sc2mac_wt_mask_9),
    .io_sc2mac_wt_mask_10(u_rt_in_io_sc2mac_wt_mask_10),
    .io_sc2mac_wt_mask_11(u_rt_in_io_sc2mac_wt_mask_11),
    .io_sc2mac_wt_mask_12(u_rt_in_io_sc2mac_wt_mask_12),
    .io_sc2mac_wt_mask_13(u_rt_in_io_sc2mac_wt_mask_13),
    .io_sc2mac_wt_mask_14(u_rt_in_io_sc2mac_wt_mask_14),
    .io_sc2mac_wt_mask_15(u_rt_in_io_sc2mac_wt_mask_15),
    .io_sc2mac_wt_mask_16(u_rt_in_io_sc2mac_wt_mask_16),
    .io_sc2mac_wt_mask_17(u_rt_in_io_sc2mac_wt_mask_17),
    .io_sc2mac_wt_mask_18(u_rt_in_io_sc2mac_wt_mask_18),
    .io_sc2mac_wt_mask_19(u_rt_in_io_sc2mac_wt_mask_19),
    .io_sc2mac_wt_mask_20(u_rt_in_io_sc2mac_wt_mask_20),
    .io_sc2mac_wt_mask_21(u_rt_in_io_sc2mac_wt_mask_21),
    .io_sc2mac_wt_mask_22(u_rt_in_io_sc2mac_wt_mask_22),
    .io_sc2mac_wt_mask_23(u_rt_in_io_sc2mac_wt_mask_23),
    .io_sc2mac_wt_mask_24(u_rt_in_io_sc2mac_wt_mask_24),
    .io_sc2mac_wt_mask_25(u_rt_in_io_sc2mac_wt_mask_25),
    .io_sc2mac_wt_mask_26(u_rt_in_io_sc2mac_wt_mask_26),
    .io_sc2mac_wt_mask_27(u_rt_in_io_sc2mac_wt_mask_27),
    .io_sc2mac_wt_mask_28(u_rt_in_io_sc2mac_wt_mask_28),
    .io_sc2mac_wt_mask_29(u_rt_in_io_sc2mac_wt_mask_29),
    .io_sc2mac_wt_mask_30(u_rt_in_io_sc2mac_wt_mask_30),
    .io_sc2mac_wt_mask_31(u_rt_in_io_sc2mac_wt_mask_31),
    .io_sc2mac_wt_mask_32(u_rt_in_io_sc2mac_wt_mask_32),
    .io_sc2mac_wt_mask_33(u_rt_in_io_sc2mac_wt_mask_33),
    .io_sc2mac_wt_mask_34(u_rt_in_io_sc2mac_wt_mask_34),
    .io_sc2mac_wt_mask_35(u_rt_in_io_sc2mac_wt_mask_35),
    .io_sc2mac_wt_mask_36(u_rt_in_io_sc2mac_wt_mask_36),
    .io_sc2mac_wt_mask_37(u_rt_in_io_sc2mac_wt_mask_37),
    .io_sc2mac_wt_mask_38(u_rt_in_io_sc2mac_wt_mask_38),
    .io_sc2mac_wt_mask_39(u_rt_in_io_sc2mac_wt_mask_39),
    .io_sc2mac_wt_mask_40(u_rt_in_io_sc2mac_wt_mask_40),
    .io_sc2mac_wt_mask_41(u_rt_in_io_sc2mac_wt_mask_41),
    .io_sc2mac_wt_mask_42(u_rt_in_io_sc2mac_wt_mask_42),
    .io_sc2mac_wt_mask_43(u_rt_in_io_sc2mac_wt_mask_43),
    .io_sc2mac_wt_mask_44(u_rt_in_io_sc2mac_wt_mask_44),
    .io_sc2mac_wt_mask_45(u_rt_in_io_sc2mac_wt_mask_45),
    .io_sc2mac_wt_mask_46(u_rt_in_io_sc2mac_wt_mask_46),
    .io_sc2mac_wt_mask_47(u_rt_in_io_sc2mac_wt_mask_47),
    .io_sc2mac_wt_mask_48(u_rt_in_io_sc2mac_wt_mask_48),
    .io_sc2mac_wt_mask_49(u_rt_in_io_sc2mac_wt_mask_49),
    .io_sc2mac_wt_mask_50(u_rt_in_io_sc2mac_wt_mask_50),
    .io_sc2mac_wt_mask_51(u_rt_in_io_sc2mac_wt_mask_51),
    .io_sc2mac_wt_mask_52(u_rt_in_io_sc2mac_wt_mask_52),
    .io_sc2mac_wt_mask_53(u_rt_in_io_sc2mac_wt_mask_53),
    .io_sc2mac_wt_mask_54(u_rt_in_io_sc2mac_wt_mask_54),
    .io_sc2mac_wt_mask_55(u_rt_in_io_sc2mac_wt_mask_55),
    .io_sc2mac_wt_mask_56(u_rt_in_io_sc2mac_wt_mask_56),
    .io_sc2mac_wt_mask_57(u_rt_in_io_sc2mac_wt_mask_57),
    .io_sc2mac_wt_mask_58(u_rt_in_io_sc2mac_wt_mask_58),
    .io_sc2mac_wt_mask_59(u_rt_in_io_sc2mac_wt_mask_59),
    .io_sc2mac_wt_mask_60(u_rt_in_io_sc2mac_wt_mask_60),
    .io_sc2mac_wt_mask_61(u_rt_in_io_sc2mac_wt_mask_61),
    .io_sc2mac_wt_mask_62(u_rt_in_io_sc2mac_wt_mask_62),
    .io_sc2mac_wt_mask_63(u_rt_in_io_sc2mac_wt_mask_63),
    .io_sc2mac_wt_mask_64(u_rt_in_io_sc2mac_wt_mask_64),
    .io_sc2mac_wt_mask_65(u_rt_in_io_sc2mac_wt_mask_65),
    .io_sc2mac_wt_mask_66(u_rt_in_io_sc2mac_wt_mask_66),
    .io_sc2mac_wt_mask_67(u_rt_in_io_sc2mac_wt_mask_67),
    .io_sc2mac_wt_mask_68(u_rt_in_io_sc2mac_wt_mask_68),
    .io_sc2mac_wt_mask_69(u_rt_in_io_sc2mac_wt_mask_69),
    .io_sc2mac_wt_mask_70(u_rt_in_io_sc2mac_wt_mask_70),
    .io_sc2mac_wt_mask_71(u_rt_in_io_sc2mac_wt_mask_71),
    .io_sc2mac_wt_mask_72(u_rt_in_io_sc2mac_wt_mask_72),
    .io_sc2mac_wt_mask_73(u_rt_in_io_sc2mac_wt_mask_73),
    .io_sc2mac_wt_mask_74(u_rt_in_io_sc2mac_wt_mask_74),
    .io_sc2mac_wt_mask_75(u_rt_in_io_sc2mac_wt_mask_75),
    .io_sc2mac_wt_mask_76(u_rt_in_io_sc2mac_wt_mask_76),
    .io_sc2mac_wt_mask_77(u_rt_in_io_sc2mac_wt_mask_77),
    .io_sc2mac_wt_mask_78(u_rt_in_io_sc2mac_wt_mask_78),
    .io_sc2mac_wt_mask_79(u_rt_in_io_sc2mac_wt_mask_79),
    .io_sc2mac_wt_mask_80(u_rt_in_io_sc2mac_wt_mask_80),
    .io_sc2mac_wt_mask_81(u_rt_in_io_sc2mac_wt_mask_81),
    .io_sc2mac_wt_mask_82(u_rt_in_io_sc2mac_wt_mask_82),
    .io_sc2mac_wt_mask_83(u_rt_in_io_sc2mac_wt_mask_83),
    .io_sc2mac_wt_mask_84(u_rt_in_io_sc2mac_wt_mask_84),
    .io_sc2mac_wt_mask_85(u_rt_in_io_sc2mac_wt_mask_85),
    .io_sc2mac_wt_mask_86(u_rt_in_io_sc2mac_wt_mask_86),
    .io_sc2mac_wt_mask_87(u_rt_in_io_sc2mac_wt_mask_87),
    .io_sc2mac_wt_mask_88(u_rt_in_io_sc2mac_wt_mask_88),
    .io_sc2mac_wt_mask_89(u_rt_in_io_sc2mac_wt_mask_89),
    .io_sc2mac_wt_mask_90(u_rt_in_io_sc2mac_wt_mask_90),
    .io_sc2mac_wt_mask_91(u_rt_in_io_sc2mac_wt_mask_91),
    .io_sc2mac_wt_mask_92(u_rt_in_io_sc2mac_wt_mask_92),
    .io_sc2mac_wt_mask_93(u_rt_in_io_sc2mac_wt_mask_93),
    .io_sc2mac_wt_mask_94(u_rt_in_io_sc2mac_wt_mask_94),
    .io_sc2mac_wt_mask_95(u_rt_in_io_sc2mac_wt_mask_95),
    .io_sc2mac_wt_mask_96(u_rt_in_io_sc2mac_wt_mask_96),
    .io_sc2mac_wt_mask_97(u_rt_in_io_sc2mac_wt_mask_97),
    .io_sc2mac_wt_mask_98(u_rt_in_io_sc2mac_wt_mask_98),
    .io_sc2mac_wt_mask_99(u_rt_in_io_sc2mac_wt_mask_99),
    .io_sc2mac_wt_mask_100(u_rt_in_io_sc2mac_wt_mask_100),
    .io_sc2mac_wt_mask_101(u_rt_in_io_sc2mac_wt_mask_101),
    .io_sc2mac_wt_mask_102(u_rt_in_io_sc2mac_wt_mask_102),
    .io_sc2mac_wt_mask_103(u_rt_in_io_sc2mac_wt_mask_103),
    .io_sc2mac_wt_mask_104(u_rt_in_io_sc2mac_wt_mask_104),
    .io_sc2mac_wt_mask_105(u_rt_in_io_sc2mac_wt_mask_105),
    .io_sc2mac_wt_mask_106(u_rt_in_io_sc2mac_wt_mask_106),
    .io_sc2mac_wt_mask_107(u_rt_in_io_sc2mac_wt_mask_107),
    .io_sc2mac_wt_mask_108(u_rt_in_io_sc2mac_wt_mask_108),
    .io_sc2mac_wt_mask_109(u_rt_in_io_sc2mac_wt_mask_109),
    .io_sc2mac_wt_mask_110(u_rt_in_io_sc2mac_wt_mask_110),
    .io_sc2mac_wt_mask_111(u_rt_in_io_sc2mac_wt_mask_111),
    .io_sc2mac_wt_mask_112(u_rt_in_io_sc2mac_wt_mask_112),
    .io_sc2mac_wt_mask_113(u_rt_in_io_sc2mac_wt_mask_113),
    .io_sc2mac_wt_mask_114(u_rt_in_io_sc2mac_wt_mask_114),
    .io_sc2mac_wt_mask_115(u_rt_in_io_sc2mac_wt_mask_115),
    .io_sc2mac_wt_mask_116(u_rt_in_io_sc2mac_wt_mask_116),
    .io_sc2mac_wt_mask_117(u_rt_in_io_sc2mac_wt_mask_117),
    .io_sc2mac_wt_mask_118(u_rt_in_io_sc2mac_wt_mask_118),
    .io_sc2mac_wt_mask_119(u_rt_in_io_sc2mac_wt_mask_119),
    .io_sc2mac_wt_mask_120(u_rt_in_io_sc2mac_wt_mask_120),
    .io_sc2mac_wt_mask_121(u_rt_in_io_sc2mac_wt_mask_121),
    .io_sc2mac_wt_mask_122(u_rt_in_io_sc2mac_wt_mask_122),
    .io_sc2mac_wt_mask_123(u_rt_in_io_sc2mac_wt_mask_123),
    .io_sc2mac_wt_mask_124(u_rt_in_io_sc2mac_wt_mask_124),
    .io_sc2mac_wt_mask_125(u_rt_in_io_sc2mac_wt_mask_125),
    .io_sc2mac_wt_mask_126(u_rt_in_io_sc2mac_wt_mask_126),
    .io_sc2mac_wt_mask_127(u_rt_in_io_sc2mac_wt_mask_127),
    .io_sc2mac_wt_sel_0(u_rt_in_io_sc2mac_wt_sel_0),
    .io_sc2mac_wt_pvld(u_rt_in_io_sc2mac_wt_pvld),
    .io_in_dat_data_0(u_rt_in_io_in_dat_data_0),
    .io_in_dat_data_1(u_rt_in_io_in_dat_data_1),
    .io_in_dat_data_2(u_rt_in_io_in_dat_data_2),
    .io_in_dat_data_3(u_rt_in_io_in_dat_data_3),
    .io_in_dat_data_4(u_rt_in_io_in_dat_data_4),
    .io_in_dat_data_5(u_rt_in_io_in_dat_data_5),
    .io_in_dat_data_6(u_rt_in_io_in_dat_data_6),
    .io_in_dat_data_7(u_rt_in_io_in_dat_data_7),
    .io_in_dat_data_8(u_rt_in_io_in_dat_data_8),
    .io_in_dat_data_9(u_rt_in_io_in_dat_data_9),
    .io_in_dat_data_10(u_rt_in_io_in_dat_data_10),
    .io_in_dat_data_11(u_rt_in_io_in_dat_data_11),
    .io_in_dat_data_12(u_rt_in_io_in_dat_data_12),
    .io_in_dat_data_13(u_rt_in_io_in_dat_data_13),
    .io_in_dat_data_14(u_rt_in_io_in_dat_data_14),
    .io_in_dat_data_15(u_rt_in_io_in_dat_data_15),
    .io_in_dat_data_16(u_rt_in_io_in_dat_data_16),
    .io_in_dat_data_17(u_rt_in_io_in_dat_data_17),
    .io_in_dat_data_18(u_rt_in_io_in_dat_data_18),
    .io_in_dat_data_19(u_rt_in_io_in_dat_data_19),
    .io_in_dat_data_20(u_rt_in_io_in_dat_data_20),
    .io_in_dat_data_21(u_rt_in_io_in_dat_data_21),
    .io_in_dat_data_22(u_rt_in_io_in_dat_data_22),
    .io_in_dat_data_23(u_rt_in_io_in_dat_data_23),
    .io_in_dat_data_24(u_rt_in_io_in_dat_data_24),
    .io_in_dat_data_25(u_rt_in_io_in_dat_data_25),
    .io_in_dat_data_26(u_rt_in_io_in_dat_data_26),
    .io_in_dat_data_27(u_rt_in_io_in_dat_data_27),
    .io_in_dat_data_28(u_rt_in_io_in_dat_data_28),
    .io_in_dat_data_29(u_rt_in_io_in_dat_data_29),
    .io_in_dat_data_30(u_rt_in_io_in_dat_data_30),
    .io_in_dat_data_31(u_rt_in_io_in_dat_data_31),
    .io_in_dat_data_32(u_rt_in_io_in_dat_data_32),
    .io_in_dat_data_33(u_rt_in_io_in_dat_data_33),
    .io_in_dat_data_34(u_rt_in_io_in_dat_data_34),
    .io_in_dat_data_35(u_rt_in_io_in_dat_data_35),
    .io_in_dat_data_36(u_rt_in_io_in_dat_data_36),
    .io_in_dat_data_37(u_rt_in_io_in_dat_data_37),
    .io_in_dat_data_38(u_rt_in_io_in_dat_data_38),
    .io_in_dat_data_39(u_rt_in_io_in_dat_data_39),
    .io_in_dat_data_40(u_rt_in_io_in_dat_data_40),
    .io_in_dat_data_41(u_rt_in_io_in_dat_data_41),
    .io_in_dat_data_42(u_rt_in_io_in_dat_data_42),
    .io_in_dat_data_43(u_rt_in_io_in_dat_data_43),
    .io_in_dat_data_44(u_rt_in_io_in_dat_data_44),
    .io_in_dat_data_45(u_rt_in_io_in_dat_data_45),
    .io_in_dat_data_46(u_rt_in_io_in_dat_data_46),
    .io_in_dat_data_47(u_rt_in_io_in_dat_data_47),
    .io_in_dat_data_48(u_rt_in_io_in_dat_data_48),
    .io_in_dat_data_49(u_rt_in_io_in_dat_data_49),
    .io_in_dat_data_50(u_rt_in_io_in_dat_data_50),
    .io_in_dat_data_51(u_rt_in_io_in_dat_data_51),
    .io_in_dat_data_52(u_rt_in_io_in_dat_data_52),
    .io_in_dat_data_53(u_rt_in_io_in_dat_data_53),
    .io_in_dat_data_54(u_rt_in_io_in_dat_data_54),
    .io_in_dat_data_55(u_rt_in_io_in_dat_data_55),
    .io_in_dat_data_56(u_rt_in_io_in_dat_data_56),
    .io_in_dat_data_57(u_rt_in_io_in_dat_data_57),
    .io_in_dat_data_58(u_rt_in_io_in_dat_data_58),
    .io_in_dat_data_59(u_rt_in_io_in_dat_data_59),
    .io_in_dat_data_60(u_rt_in_io_in_dat_data_60),
    .io_in_dat_data_61(u_rt_in_io_in_dat_data_61),
    .io_in_dat_data_62(u_rt_in_io_in_dat_data_62),
    .io_in_dat_data_63(u_rt_in_io_in_dat_data_63),
    .io_in_dat_data_64(u_rt_in_io_in_dat_data_64),
    .io_in_dat_data_65(u_rt_in_io_in_dat_data_65),
    .io_in_dat_data_66(u_rt_in_io_in_dat_data_66),
    .io_in_dat_data_67(u_rt_in_io_in_dat_data_67),
    .io_in_dat_data_68(u_rt_in_io_in_dat_data_68),
    .io_in_dat_data_69(u_rt_in_io_in_dat_data_69),
    .io_in_dat_data_70(u_rt_in_io_in_dat_data_70),
    .io_in_dat_data_71(u_rt_in_io_in_dat_data_71),
    .io_in_dat_data_72(u_rt_in_io_in_dat_data_72),
    .io_in_dat_data_73(u_rt_in_io_in_dat_data_73),
    .io_in_dat_data_74(u_rt_in_io_in_dat_data_74),
    .io_in_dat_data_75(u_rt_in_io_in_dat_data_75),
    .io_in_dat_data_76(u_rt_in_io_in_dat_data_76),
    .io_in_dat_data_77(u_rt_in_io_in_dat_data_77),
    .io_in_dat_data_78(u_rt_in_io_in_dat_data_78),
    .io_in_dat_data_79(u_rt_in_io_in_dat_data_79),
    .io_in_dat_data_80(u_rt_in_io_in_dat_data_80),
    .io_in_dat_data_81(u_rt_in_io_in_dat_data_81),
    .io_in_dat_data_82(u_rt_in_io_in_dat_data_82),
    .io_in_dat_data_83(u_rt_in_io_in_dat_data_83),
    .io_in_dat_data_84(u_rt_in_io_in_dat_data_84),
    .io_in_dat_data_85(u_rt_in_io_in_dat_data_85),
    .io_in_dat_data_86(u_rt_in_io_in_dat_data_86),
    .io_in_dat_data_87(u_rt_in_io_in_dat_data_87),
    .io_in_dat_data_88(u_rt_in_io_in_dat_data_88),
    .io_in_dat_data_89(u_rt_in_io_in_dat_data_89),
    .io_in_dat_data_90(u_rt_in_io_in_dat_data_90),
    .io_in_dat_data_91(u_rt_in_io_in_dat_data_91),
    .io_in_dat_data_92(u_rt_in_io_in_dat_data_92),
    .io_in_dat_data_93(u_rt_in_io_in_dat_data_93),
    .io_in_dat_data_94(u_rt_in_io_in_dat_data_94),
    .io_in_dat_data_95(u_rt_in_io_in_dat_data_95),
    .io_in_dat_data_96(u_rt_in_io_in_dat_data_96),
    .io_in_dat_data_97(u_rt_in_io_in_dat_data_97),
    .io_in_dat_data_98(u_rt_in_io_in_dat_data_98),
    .io_in_dat_data_99(u_rt_in_io_in_dat_data_99),
    .io_in_dat_data_100(u_rt_in_io_in_dat_data_100),
    .io_in_dat_data_101(u_rt_in_io_in_dat_data_101),
    .io_in_dat_data_102(u_rt_in_io_in_dat_data_102),
    .io_in_dat_data_103(u_rt_in_io_in_dat_data_103),
    .io_in_dat_data_104(u_rt_in_io_in_dat_data_104),
    .io_in_dat_data_105(u_rt_in_io_in_dat_data_105),
    .io_in_dat_data_106(u_rt_in_io_in_dat_data_106),
    .io_in_dat_data_107(u_rt_in_io_in_dat_data_107),
    .io_in_dat_data_108(u_rt_in_io_in_dat_data_108),
    .io_in_dat_data_109(u_rt_in_io_in_dat_data_109),
    .io_in_dat_data_110(u_rt_in_io_in_dat_data_110),
    .io_in_dat_data_111(u_rt_in_io_in_dat_data_111),
    .io_in_dat_data_112(u_rt_in_io_in_dat_data_112),
    .io_in_dat_data_113(u_rt_in_io_in_dat_data_113),
    .io_in_dat_data_114(u_rt_in_io_in_dat_data_114),
    .io_in_dat_data_115(u_rt_in_io_in_dat_data_115),
    .io_in_dat_data_116(u_rt_in_io_in_dat_data_116),
    .io_in_dat_data_117(u_rt_in_io_in_dat_data_117),
    .io_in_dat_data_118(u_rt_in_io_in_dat_data_118),
    .io_in_dat_data_119(u_rt_in_io_in_dat_data_119),
    .io_in_dat_data_120(u_rt_in_io_in_dat_data_120),
    .io_in_dat_data_121(u_rt_in_io_in_dat_data_121),
    .io_in_dat_data_122(u_rt_in_io_in_dat_data_122),
    .io_in_dat_data_123(u_rt_in_io_in_dat_data_123),
    .io_in_dat_data_124(u_rt_in_io_in_dat_data_124),
    .io_in_dat_data_125(u_rt_in_io_in_dat_data_125),
    .io_in_dat_data_126(u_rt_in_io_in_dat_data_126),
    .io_in_dat_data_127(u_rt_in_io_in_dat_data_127),
    .io_in_dat_mask_0(u_rt_in_io_in_dat_mask_0),
    .io_in_dat_mask_1(u_rt_in_io_in_dat_mask_1),
    .io_in_dat_mask_2(u_rt_in_io_in_dat_mask_2),
    .io_in_dat_mask_3(u_rt_in_io_in_dat_mask_3),
    .io_in_dat_mask_4(u_rt_in_io_in_dat_mask_4),
    .io_in_dat_mask_5(u_rt_in_io_in_dat_mask_5),
    .io_in_dat_mask_6(u_rt_in_io_in_dat_mask_6),
    .io_in_dat_mask_7(u_rt_in_io_in_dat_mask_7),
    .io_in_dat_mask_8(u_rt_in_io_in_dat_mask_8),
    .io_in_dat_mask_9(u_rt_in_io_in_dat_mask_9),
    .io_in_dat_mask_10(u_rt_in_io_in_dat_mask_10),
    .io_in_dat_mask_11(u_rt_in_io_in_dat_mask_11),
    .io_in_dat_mask_12(u_rt_in_io_in_dat_mask_12),
    .io_in_dat_mask_13(u_rt_in_io_in_dat_mask_13),
    .io_in_dat_mask_14(u_rt_in_io_in_dat_mask_14),
    .io_in_dat_mask_15(u_rt_in_io_in_dat_mask_15),
    .io_in_dat_mask_16(u_rt_in_io_in_dat_mask_16),
    .io_in_dat_mask_17(u_rt_in_io_in_dat_mask_17),
    .io_in_dat_mask_18(u_rt_in_io_in_dat_mask_18),
    .io_in_dat_mask_19(u_rt_in_io_in_dat_mask_19),
    .io_in_dat_mask_20(u_rt_in_io_in_dat_mask_20),
    .io_in_dat_mask_21(u_rt_in_io_in_dat_mask_21),
    .io_in_dat_mask_22(u_rt_in_io_in_dat_mask_22),
    .io_in_dat_mask_23(u_rt_in_io_in_dat_mask_23),
    .io_in_dat_mask_24(u_rt_in_io_in_dat_mask_24),
    .io_in_dat_mask_25(u_rt_in_io_in_dat_mask_25),
    .io_in_dat_mask_26(u_rt_in_io_in_dat_mask_26),
    .io_in_dat_mask_27(u_rt_in_io_in_dat_mask_27),
    .io_in_dat_mask_28(u_rt_in_io_in_dat_mask_28),
    .io_in_dat_mask_29(u_rt_in_io_in_dat_mask_29),
    .io_in_dat_mask_30(u_rt_in_io_in_dat_mask_30),
    .io_in_dat_mask_31(u_rt_in_io_in_dat_mask_31),
    .io_in_dat_mask_32(u_rt_in_io_in_dat_mask_32),
    .io_in_dat_mask_33(u_rt_in_io_in_dat_mask_33),
    .io_in_dat_mask_34(u_rt_in_io_in_dat_mask_34),
    .io_in_dat_mask_35(u_rt_in_io_in_dat_mask_35),
    .io_in_dat_mask_36(u_rt_in_io_in_dat_mask_36),
    .io_in_dat_mask_37(u_rt_in_io_in_dat_mask_37),
    .io_in_dat_mask_38(u_rt_in_io_in_dat_mask_38),
    .io_in_dat_mask_39(u_rt_in_io_in_dat_mask_39),
    .io_in_dat_mask_40(u_rt_in_io_in_dat_mask_40),
    .io_in_dat_mask_41(u_rt_in_io_in_dat_mask_41),
    .io_in_dat_mask_42(u_rt_in_io_in_dat_mask_42),
    .io_in_dat_mask_43(u_rt_in_io_in_dat_mask_43),
    .io_in_dat_mask_44(u_rt_in_io_in_dat_mask_44),
    .io_in_dat_mask_45(u_rt_in_io_in_dat_mask_45),
    .io_in_dat_mask_46(u_rt_in_io_in_dat_mask_46),
    .io_in_dat_mask_47(u_rt_in_io_in_dat_mask_47),
    .io_in_dat_mask_48(u_rt_in_io_in_dat_mask_48),
    .io_in_dat_mask_49(u_rt_in_io_in_dat_mask_49),
    .io_in_dat_mask_50(u_rt_in_io_in_dat_mask_50),
    .io_in_dat_mask_51(u_rt_in_io_in_dat_mask_51),
    .io_in_dat_mask_52(u_rt_in_io_in_dat_mask_52),
    .io_in_dat_mask_53(u_rt_in_io_in_dat_mask_53),
    .io_in_dat_mask_54(u_rt_in_io_in_dat_mask_54),
    .io_in_dat_mask_55(u_rt_in_io_in_dat_mask_55),
    .io_in_dat_mask_56(u_rt_in_io_in_dat_mask_56),
    .io_in_dat_mask_57(u_rt_in_io_in_dat_mask_57),
    .io_in_dat_mask_58(u_rt_in_io_in_dat_mask_58),
    .io_in_dat_mask_59(u_rt_in_io_in_dat_mask_59),
    .io_in_dat_mask_60(u_rt_in_io_in_dat_mask_60),
    .io_in_dat_mask_61(u_rt_in_io_in_dat_mask_61),
    .io_in_dat_mask_62(u_rt_in_io_in_dat_mask_62),
    .io_in_dat_mask_63(u_rt_in_io_in_dat_mask_63),
    .io_in_dat_mask_64(u_rt_in_io_in_dat_mask_64),
    .io_in_dat_mask_65(u_rt_in_io_in_dat_mask_65),
    .io_in_dat_mask_66(u_rt_in_io_in_dat_mask_66),
    .io_in_dat_mask_67(u_rt_in_io_in_dat_mask_67),
    .io_in_dat_mask_68(u_rt_in_io_in_dat_mask_68),
    .io_in_dat_mask_69(u_rt_in_io_in_dat_mask_69),
    .io_in_dat_mask_70(u_rt_in_io_in_dat_mask_70),
    .io_in_dat_mask_71(u_rt_in_io_in_dat_mask_71),
    .io_in_dat_mask_72(u_rt_in_io_in_dat_mask_72),
    .io_in_dat_mask_73(u_rt_in_io_in_dat_mask_73),
    .io_in_dat_mask_74(u_rt_in_io_in_dat_mask_74),
    .io_in_dat_mask_75(u_rt_in_io_in_dat_mask_75),
    .io_in_dat_mask_76(u_rt_in_io_in_dat_mask_76),
    .io_in_dat_mask_77(u_rt_in_io_in_dat_mask_77),
    .io_in_dat_mask_78(u_rt_in_io_in_dat_mask_78),
    .io_in_dat_mask_79(u_rt_in_io_in_dat_mask_79),
    .io_in_dat_mask_80(u_rt_in_io_in_dat_mask_80),
    .io_in_dat_mask_81(u_rt_in_io_in_dat_mask_81),
    .io_in_dat_mask_82(u_rt_in_io_in_dat_mask_82),
    .io_in_dat_mask_83(u_rt_in_io_in_dat_mask_83),
    .io_in_dat_mask_84(u_rt_in_io_in_dat_mask_84),
    .io_in_dat_mask_85(u_rt_in_io_in_dat_mask_85),
    .io_in_dat_mask_86(u_rt_in_io_in_dat_mask_86),
    .io_in_dat_mask_87(u_rt_in_io_in_dat_mask_87),
    .io_in_dat_mask_88(u_rt_in_io_in_dat_mask_88),
    .io_in_dat_mask_89(u_rt_in_io_in_dat_mask_89),
    .io_in_dat_mask_90(u_rt_in_io_in_dat_mask_90),
    .io_in_dat_mask_91(u_rt_in_io_in_dat_mask_91),
    .io_in_dat_mask_92(u_rt_in_io_in_dat_mask_92),
    .io_in_dat_mask_93(u_rt_in_io_in_dat_mask_93),
    .io_in_dat_mask_94(u_rt_in_io_in_dat_mask_94),
    .io_in_dat_mask_95(u_rt_in_io_in_dat_mask_95),
    .io_in_dat_mask_96(u_rt_in_io_in_dat_mask_96),
    .io_in_dat_mask_97(u_rt_in_io_in_dat_mask_97),
    .io_in_dat_mask_98(u_rt_in_io_in_dat_mask_98),
    .io_in_dat_mask_99(u_rt_in_io_in_dat_mask_99),
    .io_in_dat_mask_100(u_rt_in_io_in_dat_mask_100),
    .io_in_dat_mask_101(u_rt_in_io_in_dat_mask_101),
    .io_in_dat_mask_102(u_rt_in_io_in_dat_mask_102),
    .io_in_dat_mask_103(u_rt_in_io_in_dat_mask_103),
    .io_in_dat_mask_104(u_rt_in_io_in_dat_mask_104),
    .io_in_dat_mask_105(u_rt_in_io_in_dat_mask_105),
    .io_in_dat_mask_106(u_rt_in_io_in_dat_mask_106),
    .io_in_dat_mask_107(u_rt_in_io_in_dat_mask_107),
    .io_in_dat_mask_108(u_rt_in_io_in_dat_mask_108),
    .io_in_dat_mask_109(u_rt_in_io_in_dat_mask_109),
    .io_in_dat_mask_110(u_rt_in_io_in_dat_mask_110),
    .io_in_dat_mask_111(u_rt_in_io_in_dat_mask_111),
    .io_in_dat_mask_112(u_rt_in_io_in_dat_mask_112),
    .io_in_dat_mask_113(u_rt_in_io_in_dat_mask_113),
    .io_in_dat_mask_114(u_rt_in_io_in_dat_mask_114),
    .io_in_dat_mask_115(u_rt_in_io_in_dat_mask_115),
    .io_in_dat_mask_116(u_rt_in_io_in_dat_mask_116),
    .io_in_dat_mask_117(u_rt_in_io_in_dat_mask_117),
    .io_in_dat_mask_118(u_rt_in_io_in_dat_mask_118),
    .io_in_dat_mask_119(u_rt_in_io_in_dat_mask_119),
    .io_in_dat_mask_120(u_rt_in_io_in_dat_mask_120),
    .io_in_dat_mask_121(u_rt_in_io_in_dat_mask_121),
    .io_in_dat_mask_122(u_rt_in_io_in_dat_mask_122),
    .io_in_dat_mask_123(u_rt_in_io_in_dat_mask_123),
    .io_in_dat_mask_124(u_rt_in_io_in_dat_mask_124),
    .io_in_dat_mask_125(u_rt_in_io_in_dat_mask_125),
    .io_in_dat_mask_126(u_rt_in_io_in_dat_mask_126),
    .io_in_dat_mask_127(u_rt_in_io_in_dat_mask_127),
    .io_in_dat_pd(u_rt_in_io_in_dat_pd),
    .io_in_dat_pvld(u_rt_in_io_in_dat_pvld),
    .io_in_dat_stripe_st(u_rt_in_io_in_dat_stripe_st),
    .io_in_dat_stripe_end(u_rt_in_io_in_dat_stripe_end),
    .io_in_wt_data_0(u_rt_in_io_in_wt_data_0),
    .io_in_wt_data_1(u_rt_in_io_in_wt_data_1),
    .io_in_wt_data_2(u_rt_in_io_in_wt_data_2),
    .io_in_wt_data_3(u_rt_in_io_in_wt_data_3),
    .io_in_wt_data_4(u_rt_in_io_in_wt_data_4),
    .io_in_wt_data_5(u_rt_in_io_in_wt_data_5),
    .io_in_wt_data_6(u_rt_in_io_in_wt_data_6),
    .io_in_wt_data_7(u_rt_in_io_in_wt_data_7),
    .io_in_wt_data_8(u_rt_in_io_in_wt_data_8),
    .io_in_wt_data_9(u_rt_in_io_in_wt_data_9),
    .io_in_wt_data_10(u_rt_in_io_in_wt_data_10),
    .io_in_wt_data_11(u_rt_in_io_in_wt_data_11),
    .io_in_wt_data_12(u_rt_in_io_in_wt_data_12),
    .io_in_wt_data_13(u_rt_in_io_in_wt_data_13),
    .io_in_wt_data_14(u_rt_in_io_in_wt_data_14),
    .io_in_wt_data_15(u_rt_in_io_in_wt_data_15),
    .io_in_wt_data_16(u_rt_in_io_in_wt_data_16),
    .io_in_wt_data_17(u_rt_in_io_in_wt_data_17),
    .io_in_wt_data_18(u_rt_in_io_in_wt_data_18),
    .io_in_wt_data_19(u_rt_in_io_in_wt_data_19),
    .io_in_wt_data_20(u_rt_in_io_in_wt_data_20),
    .io_in_wt_data_21(u_rt_in_io_in_wt_data_21),
    .io_in_wt_data_22(u_rt_in_io_in_wt_data_22),
    .io_in_wt_data_23(u_rt_in_io_in_wt_data_23),
    .io_in_wt_data_24(u_rt_in_io_in_wt_data_24),
    .io_in_wt_data_25(u_rt_in_io_in_wt_data_25),
    .io_in_wt_data_26(u_rt_in_io_in_wt_data_26),
    .io_in_wt_data_27(u_rt_in_io_in_wt_data_27),
    .io_in_wt_data_28(u_rt_in_io_in_wt_data_28),
    .io_in_wt_data_29(u_rt_in_io_in_wt_data_29),
    .io_in_wt_data_30(u_rt_in_io_in_wt_data_30),
    .io_in_wt_data_31(u_rt_in_io_in_wt_data_31),
    .io_in_wt_data_32(u_rt_in_io_in_wt_data_32),
    .io_in_wt_data_33(u_rt_in_io_in_wt_data_33),
    .io_in_wt_data_34(u_rt_in_io_in_wt_data_34),
    .io_in_wt_data_35(u_rt_in_io_in_wt_data_35),
    .io_in_wt_data_36(u_rt_in_io_in_wt_data_36),
    .io_in_wt_data_37(u_rt_in_io_in_wt_data_37),
    .io_in_wt_data_38(u_rt_in_io_in_wt_data_38),
    .io_in_wt_data_39(u_rt_in_io_in_wt_data_39),
    .io_in_wt_data_40(u_rt_in_io_in_wt_data_40),
    .io_in_wt_data_41(u_rt_in_io_in_wt_data_41),
    .io_in_wt_data_42(u_rt_in_io_in_wt_data_42),
    .io_in_wt_data_43(u_rt_in_io_in_wt_data_43),
    .io_in_wt_data_44(u_rt_in_io_in_wt_data_44),
    .io_in_wt_data_45(u_rt_in_io_in_wt_data_45),
    .io_in_wt_data_46(u_rt_in_io_in_wt_data_46),
    .io_in_wt_data_47(u_rt_in_io_in_wt_data_47),
    .io_in_wt_data_48(u_rt_in_io_in_wt_data_48),
    .io_in_wt_data_49(u_rt_in_io_in_wt_data_49),
    .io_in_wt_data_50(u_rt_in_io_in_wt_data_50),
    .io_in_wt_data_51(u_rt_in_io_in_wt_data_51),
    .io_in_wt_data_52(u_rt_in_io_in_wt_data_52),
    .io_in_wt_data_53(u_rt_in_io_in_wt_data_53),
    .io_in_wt_data_54(u_rt_in_io_in_wt_data_54),
    .io_in_wt_data_55(u_rt_in_io_in_wt_data_55),
    .io_in_wt_data_56(u_rt_in_io_in_wt_data_56),
    .io_in_wt_data_57(u_rt_in_io_in_wt_data_57),
    .io_in_wt_data_58(u_rt_in_io_in_wt_data_58),
    .io_in_wt_data_59(u_rt_in_io_in_wt_data_59),
    .io_in_wt_data_60(u_rt_in_io_in_wt_data_60),
    .io_in_wt_data_61(u_rt_in_io_in_wt_data_61),
    .io_in_wt_data_62(u_rt_in_io_in_wt_data_62),
    .io_in_wt_data_63(u_rt_in_io_in_wt_data_63),
    .io_in_wt_data_64(u_rt_in_io_in_wt_data_64),
    .io_in_wt_data_65(u_rt_in_io_in_wt_data_65),
    .io_in_wt_data_66(u_rt_in_io_in_wt_data_66),
    .io_in_wt_data_67(u_rt_in_io_in_wt_data_67),
    .io_in_wt_data_68(u_rt_in_io_in_wt_data_68),
    .io_in_wt_data_69(u_rt_in_io_in_wt_data_69),
    .io_in_wt_data_70(u_rt_in_io_in_wt_data_70),
    .io_in_wt_data_71(u_rt_in_io_in_wt_data_71),
    .io_in_wt_data_72(u_rt_in_io_in_wt_data_72),
    .io_in_wt_data_73(u_rt_in_io_in_wt_data_73),
    .io_in_wt_data_74(u_rt_in_io_in_wt_data_74),
    .io_in_wt_data_75(u_rt_in_io_in_wt_data_75),
    .io_in_wt_data_76(u_rt_in_io_in_wt_data_76),
    .io_in_wt_data_77(u_rt_in_io_in_wt_data_77),
    .io_in_wt_data_78(u_rt_in_io_in_wt_data_78),
    .io_in_wt_data_79(u_rt_in_io_in_wt_data_79),
    .io_in_wt_data_80(u_rt_in_io_in_wt_data_80),
    .io_in_wt_data_81(u_rt_in_io_in_wt_data_81),
    .io_in_wt_data_82(u_rt_in_io_in_wt_data_82),
    .io_in_wt_data_83(u_rt_in_io_in_wt_data_83),
    .io_in_wt_data_84(u_rt_in_io_in_wt_data_84),
    .io_in_wt_data_85(u_rt_in_io_in_wt_data_85),
    .io_in_wt_data_86(u_rt_in_io_in_wt_data_86),
    .io_in_wt_data_87(u_rt_in_io_in_wt_data_87),
    .io_in_wt_data_88(u_rt_in_io_in_wt_data_88),
    .io_in_wt_data_89(u_rt_in_io_in_wt_data_89),
    .io_in_wt_data_90(u_rt_in_io_in_wt_data_90),
    .io_in_wt_data_91(u_rt_in_io_in_wt_data_91),
    .io_in_wt_data_92(u_rt_in_io_in_wt_data_92),
    .io_in_wt_data_93(u_rt_in_io_in_wt_data_93),
    .io_in_wt_data_94(u_rt_in_io_in_wt_data_94),
    .io_in_wt_data_95(u_rt_in_io_in_wt_data_95),
    .io_in_wt_data_96(u_rt_in_io_in_wt_data_96),
    .io_in_wt_data_97(u_rt_in_io_in_wt_data_97),
    .io_in_wt_data_98(u_rt_in_io_in_wt_data_98),
    .io_in_wt_data_99(u_rt_in_io_in_wt_data_99),
    .io_in_wt_data_100(u_rt_in_io_in_wt_data_100),
    .io_in_wt_data_101(u_rt_in_io_in_wt_data_101),
    .io_in_wt_data_102(u_rt_in_io_in_wt_data_102),
    .io_in_wt_data_103(u_rt_in_io_in_wt_data_103),
    .io_in_wt_data_104(u_rt_in_io_in_wt_data_104),
    .io_in_wt_data_105(u_rt_in_io_in_wt_data_105),
    .io_in_wt_data_106(u_rt_in_io_in_wt_data_106),
    .io_in_wt_data_107(u_rt_in_io_in_wt_data_107),
    .io_in_wt_data_108(u_rt_in_io_in_wt_data_108),
    .io_in_wt_data_109(u_rt_in_io_in_wt_data_109),
    .io_in_wt_data_110(u_rt_in_io_in_wt_data_110),
    .io_in_wt_data_111(u_rt_in_io_in_wt_data_111),
    .io_in_wt_data_112(u_rt_in_io_in_wt_data_112),
    .io_in_wt_data_113(u_rt_in_io_in_wt_data_113),
    .io_in_wt_data_114(u_rt_in_io_in_wt_data_114),
    .io_in_wt_data_115(u_rt_in_io_in_wt_data_115),
    .io_in_wt_data_116(u_rt_in_io_in_wt_data_116),
    .io_in_wt_data_117(u_rt_in_io_in_wt_data_117),
    .io_in_wt_data_118(u_rt_in_io_in_wt_data_118),
    .io_in_wt_data_119(u_rt_in_io_in_wt_data_119),
    .io_in_wt_data_120(u_rt_in_io_in_wt_data_120),
    .io_in_wt_data_121(u_rt_in_io_in_wt_data_121),
    .io_in_wt_data_122(u_rt_in_io_in_wt_data_122),
    .io_in_wt_data_123(u_rt_in_io_in_wt_data_123),
    .io_in_wt_data_124(u_rt_in_io_in_wt_data_124),
    .io_in_wt_data_125(u_rt_in_io_in_wt_data_125),
    .io_in_wt_data_126(u_rt_in_io_in_wt_data_126),
    .io_in_wt_data_127(u_rt_in_io_in_wt_data_127),
    .io_in_wt_mask_0(u_rt_in_io_in_wt_mask_0),
    .io_in_wt_mask_1(u_rt_in_io_in_wt_mask_1),
    .io_in_wt_mask_2(u_rt_in_io_in_wt_mask_2),
    .io_in_wt_mask_3(u_rt_in_io_in_wt_mask_3),
    .io_in_wt_mask_4(u_rt_in_io_in_wt_mask_4),
    .io_in_wt_mask_5(u_rt_in_io_in_wt_mask_5),
    .io_in_wt_mask_6(u_rt_in_io_in_wt_mask_6),
    .io_in_wt_mask_7(u_rt_in_io_in_wt_mask_7),
    .io_in_wt_mask_8(u_rt_in_io_in_wt_mask_8),
    .io_in_wt_mask_9(u_rt_in_io_in_wt_mask_9),
    .io_in_wt_mask_10(u_rt_in_io_in_wt_mask_10),
    .io_in_wt_mask_11(u_rt_in_io_in_wt_mask_11),
    .io_in_wt_mask_12(u_rt_in_io_in_wt_mask_12),
    .io_in_wt_mask_13(u_rt_in_io_in_wt_mask_13),
    .io_in_wt_mask_14(u_rt_in_io_in_wt_mask_14),
    .io_in_wt_mask_15(u_rt_in_io_in_wt_mask_15),
    .io_in_wt_mask_16(u_rt_in_io_in_wt_mask_16),
    .io_in_wt_mask_17(u_rt_in_io_in_wt_mask_17),
    .io_in_wt_mask_18(u_rt_in_io_in_wt_mask_18),
    .io_in_wt_mask_19(u_rt_in_io_in_wt_mask_19),
    .io_in_wt_mask_20(u_rt_in_io_in_wt_mask_20),
    .io_in_wt_mask_21(u_rt_in_io_in_wt_mask_21),
    .io_in_wt_mask_22(u_rt_in_io_in_wt_mask_22),
    .io_in_wt_mask_23(u_rt_in_io_in_wt_mask_23),
    .io_in_wt_mask_24(u_rt_in_io_in_wt_mask_24),
    .io_in_wt_mask_25(u_rt_in_io_in_wt_mask_25),
    .io_in_wt_mask_26(u_rt_in_io_in_wt_mask_26),
    .io_in_wt_mask_27(u_rt_in_io_in_wt_mask_27),
    .io_in_wt_mask_28(u_rt_in_io_in_wt_mask_28),
    .io_in_wt_mask_29(u_rt_in_io_in_wt_mask_29),
    .io_in_wt_mask_30(u_rt_in_io_in_wt_mask_30),
    .io_in_wt_mask_31(u_rt_in_io_in_wt_mask_31),
    .io_in_wt_mask_32(u_rt_in_io_in_wt_mask_32),
    .io_in_wt_mask_33(u_rt_in_io_in_wt_mask_33),
    .io_in_wt_mask_34(u_rt_in_io_in_wt_mask_34),
    .io_in_wt_mask_35(u_rt_in_io_in_wt_mask_35),
    .io_in_wt_mask_36(u_rt_in_io_in_wt_mask_36),
    .io_in_wt_mask_37(u_rt_in_io_in_wt_mask_37),
    .io_in_wt_mask_38(u_rt_in_io_in_wt_mask_38),
    .io_in_wt_mask_39(u_rt_in_io_in_wt_mask_39),
    .io_in_wt_mask_40(u_rt_in_io_in_wt_mask_40),
    .io_in_wt_mask_41(u_rt_in_io_in_wt_mask_41),
    .io_in_wt_mask_42(u_rt_in_io_in_wt_mask_42),
    .io_in_wt_mask_43(u_rt_in_io_in_wt_mask_43),
    .io_in_wt_mask_44(u_rt_in_io_in_wt_mask_44),
    .io_in_wt_mask_45(u_rt_in_io_in_wt_mask_45),
    .io_in_wt_mask_46(u_rt_in_io_in_wt_mask_46),
    .io_in_wt_mask_47(u_rt_in_io_in_wt_mask_47),
    .io_in_wt_mask_48(u_rt_in_io_in_wt_mask_48),
    .io_in_wt_mask_49(u_rt_in_io_in_wt_mask_49),
    .io_in_wt_mask_50(u_rt_in_io_in_wt_mask_50),
    .io_in_wt_mask_51(u_rt_in_io_in_wt_mask_51),
    .io_in_wt_mask_52(u_rt_in_io_in_wt_mask_52),
    .io_in_wt_mask_53(u_rt_in_io_in_wt_mask_53),
    .io_in_wt_mask_54(u_rt_in_io_in_wt_mask_54),
    .io_in_wt_mask_55(u_rt_in_io_in_wt_mask_55),
    .io_in_wt_mask_56(u_rt_in_io_in_wt_mask_56),
    .io_in_wt_mask_57(u_rt_in_io_in_wt_mask_57),
    .io_in_wt_mask_58(u_rt_in_io_in_wt_mask_58),
    .io_in_wt_mask_59(u_rt_in_io_in_wt_mask_59),
    .io_in_wt_mask_60(u_rt_in_io_in_wt_mask_60),
    .io_in_wt_mask_61(u_rt_in_io_in_wt_mask_61),
    .io_in_wt_mask_62(u_rt_in_io_in_wt_mask_62),
    .io_in_wt_mask_63(u_rt_in_io_in_wt_mask_63),
    .io_in_wt_mask_64(u_rt_in_io_in_wt_mask_64),
    .io_in_wt_mask_65(u_rt_in_io_in_wt_mask_65),
    .io_in_wt_mask_66(u_rt_in_io_in_wt_mask_66),
    .io_in_wt_mask_67(u_rt_in_io_in_wt_mask_67),
    .io_in_wt_mask_68(u_rt_in_io_in_wt_mask_68),
    .io_in_wt_mask_69(u_rt_in_io_in_wt_mask_69),
    .io_in_wt_mask_70(u_rt_in_io_in_wt_mask_70),
    .io_in_wt_mask_71(u_rt_in_io_in_wt_mask_71),
    .io_in_wt_mask_72(u_rt_in_io_in_wt_mask_72),
    .io_in_wt_mask_73(u_rt_in_io_in_wt_mask_73),
    .io_in_wt_mask_74(u_rt_in_io_in_wt_mask_74),
    .io_in_wt_mask_75(u_rt_in_io_in_wt_mask_75),
    .io_in_wt_mask_76(u_rt_in_io_in_wt_mask_76),
    .io_in_wt_mask_77(u_rt_in_io_in_wt_mask_77),
    .io_in_wt_mask_78(u_rt_in_io_in_wt_mask_78),
    .io_in_wt_mask_79(u_rt_in_io_in_wt_mask_79),
    .io_in_wt_mask_80(u_rt_in_io_in_wt_mask_80),
    .io_in_wt_mask_81(u_rt_in_io_in_wt_mask_81),
    .io_in_wt_mask_82(u_rt_in_io_in_wt_mask_82),
    .io_in_wt_mask_83(u_rt_in_io_in_wt_mask_83),
    .io_in_wt_mask_84(u_rt_in_io_in_wt_mask_84),
    .io_in_wt_mask_85(u_rt_in_io_in_wt_mask_85),
    .io_in_wt_mask_86(u_rt_in_io_in_wt_mask_86),
    .io_in_wt_mask_87(u_rt_in_io_in_wt_mask_87),
    .io_in_wt_mask_88(u_rt_in_io_in_wt_mask_88),
    .io_in_wt_mask_89(u_rt_in_io_in_wt_mask_89),
    .io_in_wt_mask_90(u_rt_in_io_in_wt_mask_90),
    .io_in_wt_mask_91(u_rt_in_io_in_wt_mask_91),
    .io_in_wt_mask_92(u_rt_in_io_in_wt_mask_92),
    .io_in_wt_mask_93(u_rt_in_io_in_wt_mask_93),
    .io_in_wt_mask_94(u_rt_in_io_in_wt_mask_94),
    .io_in_wt_mask_95(u_rt_in_io_in_wt_mask_95),
    .io_in_wt_mask_96(u_rt_in_io_in_wt_mask_96),
    .io_in_wt_mask_97(u_rt_in_io_in_wt_mask_97),
    .io_in_wt_mask_98(u_rt_in_io_in_wt_mask_98),
    .io_in_wt_mask_99(u_rt_in_io_in_wt_mask_99),
    .io_in_wt_mask_100(u_rt_in_io_in_wt_mask_100),
    .io_in_wt_mask_101(u_rt_in_io_in_wt_mask_101),
    .io_in_wt_mask_102(u_rt_in_io_in_wt_mask_102),
    .io_in_wt_mask_103(u_rt_in_io_in_wt_mask_103),
    .io_in_wt_mask_104(u_rt_in_io_in_wt_mask_104),
    .io_in_wt_mask_105(u_rt_in_io_in_wt_mask_105),
    .io_in_wt_mask_106(u_rt_in_io_in_wt_mask_106),
    .io_in_wt_mask_107(u_rt_in_io_in_wt_mask_107),
    .io_in_wt_mask_108(u_rt_in_io_in_wt_mask_108),
    .io_in_wt_mask_109(u_rt_in_io_in_wt_mask_109),
    .io_in_wt_mask_110(u_rt_in_io_in_wt_mask_110),
    .io_in_wt_mask_111(u_rt_in_io_in_wt_mask_111),
    .io_in_wt_mask_112(u_rt_in_io_in_wt_mask_112),
    .io_in_wt_mask_113(u_rt_in_io_in_wt_mask_113),
    .io_in_wt_mask_114(u_rt_in_io_in_wt_mask_114),
    .io_in_wt_mask_115(u_rt_in_io_in_wt_mask_115),
    .io_in_wt_mask_116(u_rt_in_io_in_wt_mask_116),
    .io_in_wt_mask_117(u_rt_in_io_in_wt_mask_117),
    .io_in_wt_mask_118(u_rt_in_io_in_wt_mask_118),
    .io_in_wt_mask_119(u_rt_in_io_in_wt_mask_119),
    .io_in_wt_mask_120(u_rt_in_io_in_wt_mask_120),
    .io_in_wt_mask_121(u_rt_in_io_in_wt_mask_121),
    .io_in_wt_mask_122(u_rt_in_io_in_wt_mask_122),
    .io_in_wt_mask_123(u_rt_in_io_in_wt_mask_123),
    .io_in_wt_mask_124(u_rt_in_io_in_wt_mask_124),
    .io_in_wt_mask_125(u_rt_in_io_in_wt_mask_125),
    .io_in_wt_mask_126(u_rt_in_io_in_wt_mask_126),
    .io_in_wt_mask_127(u_rt_in_io_in_wt_mask_127),
    .io_in_wt_sel_0(u_rt_in_io_in_wt_sel_0),
    .io_in_wt_pvld(u_rt_in_io_in_wt_pvld)
  );
  NV_NVDLA_CMAC_CORE_active u_active ( // @[NV_NVDLA_CMAC_core.scala 82:26]
    .clock(u_active_clock),
    .reset(u_active_reset),
    .io_in_dat_data_0(u_active_io_in_dat_data_0),
    .io_in_dat_data_1(u_active_io_in_dat_data_1),
    .io_in_dat_data_2(u_active_io_in_dat_data_2),
    .io_in_dat_data_3(u_active_io_in_dat_data_3),
    .io_in_dat_data_4(u_active_io_in_dat_data_4),
    .io_in_dat_data_5(u_active_io_in_dat_data_5),
    .io_in_dat_data_6(u_active_io_in_dat_data_6),
    .io_in_dat_data_7(u_active_io_in_dat_data_7),
    .io_in_dat_data_8(u_active_io_in_dat_data_8),
    .io_in_dat_data_9(u_active_io_in_dat_data_9),
    .io_in_dat_data_10(u_active_io_in_dat_data_10),
    .io_in_dat_data_11(u_active_io_in_dat_data_11),
    .io_in_dat_data_12(u_active_io_in_dat_data_12),
    .io_in_dat_data_13(u_active_io_in_dat_data_13),
    .io_in_dat_data_14(u_active_io_in_dat_data_14),
    .io_in_dat_data_15(u_active_io_in_dat_data_15),
    .io_in_dat_data_16(u_active_io_in_dat_data_16),
    .io_in_dat_data_17(u_active_io_in_dat_data_17),
    .io_in_dat_data_18(u_active_io_in_dat_data_18),
    .io_in_dat_data_19(u_active_io_in_dat_data_19),
    .io_in_dat_data_20(u_active_io_in_dat_data_20),
    .io_in_dat_data_21(u_active_io_in_dat_data_21),
    .io_in_dat_data_22(u_active_io_in_dat_data_22),
    .io_in_dat_data_23(u_active_io_in_dat_data_23),
    .io_in_dat_data_24(u_active_io_in_dat_data_24),
    .io_in_dat_data_25(u_active_io_in_dat_data_25),
    .io_in_dat_data_26(u_active_io_in_dat_data_26),
    .io_in_dat_data_27(u_active_io_in_dat_data_27),
    .io_in_dat_data_28(u_active_io_in_dat_data_28),
    .io_in_dat_data_29(u_active_io_in_dat_data_29),
    .io_in_dat_data_30(u_active_io_in_dat_data_30),
    .io_in_dat_data_31(u_active_io_in_dat_data_31),
    .io_in_dat_data_32(u_active_io_in_dat_data_32),
    .io_in_dat_data_33(u_active_io_in_dat_data_33),
    .io_in_dat_data_34(u_active_io_in_dat_data_34),
    .io_in_dat_data_35(u_active_io_in_dat_data_35),
    .io_in_dat_data_36(u_active_io_in_dat_data_36),
    .io_in_dat_data_37(u_active_io_in_dat_data_37),
    .io_in_dat_data_38(u_active_io_in_dat_data_38),
    .io_in_dat_data_39(u_active_io_in_dat_data_39),
    .io_in_dat_data_40(u_active_io_in_dat_data_40),
    .io_in_dat_data_41(u_active_io_in_dat_data_41),
    .io_in_dat_data_42(u_active_io_in_dat_data_42),
    .io_in_dat_data_43(u_active_io_in_dat_data_43),
    .io_in_dat_data_44(u_active_io_in_dat_data_44),
    .io_in_dat_data_45(u_active_io_in_dat_data_45),
    .io_in_dat_data_46(u_active_io_in_dat_data_46),
    .io_in_dat_data_47(u_active_io_in_dat_data_47),
    .io_in_dat_data_48(u_active_io_in_dat_data_48),
    .io_in_dat_data_49(u_active_io_in_dat_data_49),
    .io_in_dat_data_50(u_active_io_in_dat_data_50),
    .io_in_dat_data_51(u_active_io_in_dat_data_51),
    .io_in_dat_data_52(u_active_io_in_dat_data_52),
    .io_in_dat_data_53(u_active_io_in_dat_data_53),
    .io_in_dat_data_54(u_active_io_in_dat_data_54),
    .io_in_dat_data_55(u_active_io_in_dat_data_55),
    .io_in_dat_data_56(u_active_io_in_dat_data_56),
    .io_in_dat_data_57(u_active_io_in_dat_data_57),
    .io_in_dat_data_58(u_active_io_in_dat_data_58),
    .io_in_dat_data_59(u_active_io_in_dat_data_59),
    .io_in_dat_data_60(u_active_io_in_dat_data_60),
    .io_in_dat_data_61(u_active_io_in_dat_data_61),
    .io_in_dat_data_62(u_active_io_in_dat_data_62),
    .io_in_dat_data_63(u_active_io_in_dat_data_63),
    .io_in_dat_data_64(u_active_io_in_dat_data_64),
    .io_in_dat_data_65(u_active_io_in_dat_data_65),
    .io_in_dat_data_66(u_active_io_in_dat_data_66),
    .io_in_dat_data_67(u_active_io_in_dat_data_67),
    .io_in_dat_data_68(u_active_io_in_dat_data_68),
    .io_in_dat_data_69(u_active_io_in_dat_data_69),
    .io_in_dat_data_70(u_active_io_in_dat_data_70),
    .io_in_dat_data_71(u_active_io_in_dat_data_71),
    .io_in_dat_data_72(u_active_io_in_dat_data_72),
    .io_in_dat_data_73(u_active_io_in_dat_data_73),
    .io_in_dat_data_74(u_active_io_in_dat_data_74),
    .io_in_dat_data_75(u_active_io_in_dat_data_75),
    .io_in_dat_data_76(u_active_io_in_dat_data_76),
    .io_in_dat_data_77(u_active_io_in_dat_data_77),
    .io_in_dat_data_78(u_active_io_in_dat_data_78),
    .io_in_dat_data_79(u_active_io_in_dat_data_79),
    .io_in_dat_data_80(u_active_io_in_dat_data_80),
    .io_in_dat_data_81(u_active_io_in_dat_data_81),
    .io_in_dat_data_82(u_active_io_in_dat_data_82),
    .io_in_dat_data_83(u_active_io_in_dat_data_83),
    .io_in_dat_data_84(u_active_io_in_dat_data_84),
    .io_in_dat_data_85(u_active_io_in_dat_data_85),
    .io_in_dat_data_86(u_active_io_in_dat_data_86),
    .io_in_dat_data_87(u_active_io_in_dat_data_87),
    .io_in_dat_data_88(u_active_io_in_dat_data_88),
    .io_in_dat_data_89(u_active_io_in_dat_data_89),
    .io_in_dat_data_90(u_active_io_in_dat_data_90),
    .io_in_dat_data_91(u_active_io_in_dat_data_91),
    .io_in_dat_data_92(u_active_io_in_dat_data_92),
    .io_in_dat_data_93(u_active_io_in_dat_data_93),
    .io_in_dat_data_94(u_active_io_in_dat_data_94),
    .io_in_dat_data_95(u_active_io_in_dat_data_95),
    .io_in_dat_data_96(u_active_io_in_dat_data_96),
    .io_in_dat_data_97(u_active_io_in_dat_data_97),
    .io_in_dat_data_98(u_active_io_in_dat_data_98),
    .io_in_dat_data_99(u_active_io_in_dat_data_99),
    .io_in_dat_data_100(u_active_io_in_dat_data_100),
    .io_in_dat_data_101(u_active_io_in_dat_data_101),
    .io_in_dat_data_102(u_active_io_in_dat_data_102),
    .io_in_dat_data_103(u_active_io_in_dat_data_103),
    .io_in_dat_data_104(u_active_io_in_dat_data_104),
    .io_in_dat_data_105(u_active_io_in_dat_data_105),
    .io_in_dat_data_106(u_active_io_in_dat_data_106),
    .io_in_dat_data_107(u_active_io_in_dat_data_107),
    .io_in_dat_data_108(u_active_io_in_dat_data_108),
    .io_in_dat_data_109(u_active_io_in_dat_data_109),
    .io_in_dat_data_110(u_active_io_in_dat_data_110),
    .io_in_dat_data_111(u_active_io_in_dat_data_111),
    .io_in_dat_data_112(u_active_io_in_dat_data_112),
    .io_in_dat_data_113(u_active_io_in_dat_data_113),
    .io_in_dat_data_114(u_active_io_in_dat_data_114),
    .io_in_dat_data_115(u_active_io_in_dat_data_115),
    .io_in_dat_data_116(u_active_io_in_dat_data_116),
    .io_in_dat_data_117(u_active_io_in_dat_data_117),
    .io_in_dat_data_118(u_active_io_in_dat_data_118),
    .io_in_dat_data_119(u_active_io_in_dat_data_119),
    .io_in_dat_data_120(u_active_io_in_dat_data_120),
    .io_in_dat_data_121(u_active_io_in_dat_data_121),
    .io_in_dat_data_122(u_active_io_in_dat_data_122),
    .io_in_dat_data_123(u_active_io_in_dat_data_123),
    .io_in_dat_data_124(u_active_io_in_dat_data_124),
    .io_in_dat_data_125(u_active_io_in_dat_data_125),
    .io_in_dat_data_126(u_active_io_in_dat_data_126),
    .io_in_dat_data_127(u_active_io_in_dat_data_127),
    .io_in_dat_mask_0(u_active_io_in_dat_mask_0),
    .io_in_dat_mask_1(u_active_io_in_dat_mask_1),
    .io_in_dat_mask_2(u_active_io_in_dat_mask_2),
    .io_in_dat_mask_3(u_active_io_in_dat_mask_3),
    .io_in_dat_mask_4(u_active_io_in_dat_mask_4),
    .io_in_dat_mask_5(u_active_io_in_dat_mask_5),
    .io_in_dat_mask_6(u_active_io_in_dat_mask_6),
    .io_in_dat_mask_7(u_active_io_in_dat_mask_7),
    .io_in_dat_mask_8(u_active_io_in_dat_mask_8),
    .io_in_dat_mask_9(u_active_io_in_dat_mask_9),
    .io_in_dat_mask_10(u_active_io_in_dat_mask_10),
    .io_in_dat_mask_11(u_active_io_in_dat_mask_11),
    .io_in_dat_mask_12(u_active_io_in_dat_mask_12),
    .io_in_dat_mask_13(u_active_io_in_dat_mask_13),
    .io_in_dat_mask_14(u_active_io_in_dat_mask_14),
    .io_in_dat_mask_15(u_active_io_in_dat_mask_15),
    .io_in_dat_mask_16(u_active_io_in_dat_mask_16),
    .io_in_dat_mask_17(u_active_io_in_dat_mask_17),
    .io_in_dat_mask_18(u_active_io_in_dat_mask_18),
    .io_in_dat_mask_19(u_active_io_in_dat_mask_19),
    .io_in_dat_mask_20(u_active_io_in_dat_mask_20),
    .io_in_dat_mask_21(u_active_io_in_dat_mask_21),
    .io_in_dat_mask_22(u_active_io_in_dat_mask_22),
    .io_in_dat_mask_23(u_active_io_in_dat_mask_23),
    .io_in_dat_mask_24(u_active_io_in_dat_mask_24),
    .io_in_dat_mask_25(u_active_io_in_dat_mask_25),
    .io_in_dat_mask_26(u_active_io_in_dat_mask_26),
    .io_in_dat_mask_27(u_active_io_in_dat_mask_27),
    .io_in_dat_mask_28(u_active_io_in_dat_mask_28),
    .io_in_dat_mask_29(u_active_io_in_dat_mask_29),
    .io_in_dat_mask_30(u_active_io_in_dat_mask_30),
    .io_in_dat_mask_31(u_active_io_in_dat_mask_31),
    .io_in_dat_mask_32(u_active_io_in_dat_mask_32),
    .io_in_dat_mask_33(u_active_io_in_dat_mask_33),
    .io_in_dat_mask_34(u_active_io_in_dat_mask_34),
    .io_in_dat_mask_35(u_active_io_in_dat_mask_35),
    .io_in_dat_mask_36(u_active_io_in_dat_mask_36),
    .io_in_dat_mask_37(u_active_io_in_dat_mask_37),
    .io_in_dat_mask_38(u_active_io_in_dat_mask_38),
    .io_in_dat_mask_39(u_active_io_in_dat_mask_39),
    .io_in_dat_mask_40(u_active_io_in_dat_mask_40),
    .io_in_dat_mask_41(u_active_io_in_dat_mask_41),
    .io_in_dat_mask_42(u_active_io_in_dat_mask_42),
    .io_in_dat_mask_43(u_active_io_in_dat_mask_43),
    .io_in_dat_mask_44(u_active_io_in_dat_mask_44),
    .io_in_dat_mask_45(u_active_io_in_dat_mask_45),
    .io_in_dat_mask_46(u_active_io_in_dat_mask_46),
    .io_in_dat_mask_47(u_active_io_in_dat_mask_47),
    .io_in_dat_mask_48(u_active_io_in_dat_mask_48),
    .io_in_dat_mask_49(u_active_io_in_dat_mask_49),
    .io_in_dat_mask_50(u_active_io_in_dat_mask_50),
    .io_in_dat_mask_51(u_active_io_in_dat_mask_51),
    .io_in_dat_mask_52(u_active_io_in_dat_mask_52),
    .io_in_dat_mask_53(u_active_io_in_dat_mask_53),
    .io_in_dat_mask_54(u_active_io_in_dat_mask_54),
    .io_in_dat_mask_55(u_active_io_in_dat_mask_55),
    .io_in_dat_mask_56(u_active_io_in_dat_mask_56),
    .io_in_dat_mask_57(u_active_io_in_dat_mask_57),
    .io_in_dat_mask_58(u_active_io_in_dat_mask_58),
    .io_in_dat_mask_59(u_active_io_in_dat_mask_59),
    .io_in_dat_mask_60(u_active_io_in_dat_mask_60),
    .io_in_dat_mask_61(u_active_io_in_dat_mask_61),
    .io_in_dat_mask_62(u_active_io_in_dat_mask_62),
    .io_in_dat_mask_63(u_active_io_in_dat_mask_63),
    .io_in_dat_mask_64(u_active_io_in_dat_mask_64),
    .io_in_dat_mask_65(u_active_io_in_dat_mask_65),
    .io_in_dat_mask_66(u_active_io_in_dat_mask_66),
    .io_in_dat_mask_67(u_active_io_in_dat_mask_67),
    .io_in_dat_mask_68(u_active_io_in_dat_mask_68),
    .io_in_dat_mask_69(u_active_io_in_dat_mask_69),
    .io_in_dat_mask_70(u_active_io_in_dat_mask_70),
    .io_in_dat_mask_71(u_active_io_in_dat_mask_71),
    .io_in_dat_mask_72(u_active_io_in_dat_mask_72),
    .io_in_dat_mask_73(u_active_io_in_dat_mask_73),
    .io_in_dat_mask_74(u_active_io_in_dat_mask_74),
    .io_in_dat_mask_75(u_active_io_in_dat_mask_75),
    .io_in_dat_mask_76(u_active_io_in_dat_mask_76),
    .io_in_dat_mask_77(u_active_io_in_dat_mask_77),
    .io_in_dat_mask_78(u_active_io_in_dat_mask_78),
    .io_in_dat_mask_79(u_active_io_in_dat_mask_79),
    .io_in_dat_mask_80(u_active_io_in_dat_mask_80),
    .io_in_dat_mask_81(u_active_io_in_dat_mask_81),
    .io_in_dat_mask_82(u_active_io_in_dat_mask_82),
    .io_in_dat_mask_83(u_active_io_in_dat_mask_83),
    .io_in_dat_mask_84(u_active_io_in_dat_mask_84),
    .io_in_dat_mask_85(u_active_io_in_dat_mask_85),
    .io_in_dat_mask_86(u_active_io_in_dat_mask_86),
    .io_in_dat_mask_87(u_active_io_in_dat_mask_87),
    .io_in_dat_mask_88(u_active_io_in_dat_mask_88),
    .io_in_dat_mask_89(u_active_io_in_dat_mask_89),
    .io_in_dat_mask_90(u_active_io_in_dat_mask_90),
    .io_in_dat_mask_91(u_active_io_in_dat_mask_91),
    .io_in_dat_mask_92(u_active_io_in_dat_mask_92),
    .io_in_dat_mask_93(u_active_io_in_dat_mask_93),
    .io_in_dat_mask_94(u_active_io_in_dat_mask_94),
    .io_in_dat_mask_95(u_active_io_in_dat_mask_95),
    .io_in_dat_mask_96(u_active_io_in_dat_mask_96),
    .io_in_dat_mask_97(u_active_io_in_dat_mask_97),
    .io_in_dat_mask_98(u_active_io_in_dat_mask_98),
    .io_in_dat_mask_99(u_active_io_in_dat_mask_99),
    .io_in_dat_mask_100(u_active_io_in_dat_mask_100),
    .io_in_dat_mask_101(u_active_io_in_dat_mask_101),
    .io_in_dat_mask_102(u_active_io_in_dat_mask_102),
    .io_in_dat_mask_103(u_active_io_in_dat_mask_103),
    .io_in_dat_mask_104(u_active_io_in_dat_mask_104),
    .io_in_dat_mask_105(u_active_io_in_dat_mask_105),
    .io_in_dat_mask_106(u_active_io_in_dat_mask_106),
    .io_in_dat_mask_107(u_active_io_in_dat_mask_107),
    .io_in_dat_mask_108(u_active_io_in_dat_mask_108),
    .io_in_dat_mask_109(u_active_io_in_dat_mask_109),
    .io_in_dat_mask_110(u_active_io_in_dat_mask_110),
    .io_in_dat_mask_111(u_active_io_in_dat_mask_111),
    .io_in_dat_mask_112(u_active_io_in_dat_mask_112),
    .io_in_dat_mask_113(u_active_io_in_dat_mask_113),
    .io_in_dat_mask_114(u_active_io_in_dat_mask_114),
    .io_in_dat_mask_115(u_active_io_in_dat_mask_115),
    .io_in_dat_mask_116(u_active_io_in_dat_mask_116),
    .io_in_dat_mask_117(u_active_io_in_dat_mask_117),
    .io_in_dat_mask_118(u_active_io_in_dat_mask_118),
    .io_in_dat_mask_119(u_active_io_in_dat_mask_119),
    .io_in_dat_mask_120(u_active_io_in_dat_mask_120),
    .io_in_dat_mask_121(u_active_io_in_dat_mask_121),
    .io_in_dat_mask_122(u_active_io_in_dat_mask_122),
    .io_in_dat_mask_123(u_active_io_in_dat_mask_123),
    .io_in_dat_mask_124(u_active_io_in_dat_mask_124),
    .io_in_dat_mask_125(u_active_io_in_dat_mask_125),
    .io_in_dat_mask_126(u_active_io_in_dat_mask_126),
    .io_in_dat_mask_127(u_active_io_in_dat_mask_127),
    .io_in_dat_pvld(u_active_io_in_dat_pvld),
    .io_in_dat_stripe_st(u_active_io_in_dat_stripe_st),
    .io_in_dat_stripe_end(u_active_io_in_dat_stripe_end),
    .io_in_wt_data_0(u_active_io_in_wt_data_0),
    .io_in_wt_data_1(u_active_io_in_wt_data_1),
    .io_in_wt_data_2(u_active_io_in_wt_data_2),
    .io_in_wt_data_3(u_active_io_in_wt_data_3),
    .io_in_wt_data_4(u_active_io_in_wt_data_4),
    .io_in_wt_data_5(u_active_io_in_wt_data_5),
    .io_in_wt_data_6(u_active_io_in_wt_data_6),
    .io_in_wt_data_7(u_active_io_in_wt_data_7),
    .io_in_wt_data_8(u_active_io_in_wt_data_8),
    .io_in_wt_data_9(u_active_io_in_wt_data_9),
    .io_in_wt_data_10(u_active_io_in_wt_data_10),
    .io_in_wt_data_11(u_active_io_in_wt_data_11),
    .io_in_wt_data_12(u_active_io_in_wt_data_12),
    .io_in_wt_data_13(u_active_io_in_wt_data_13),
    .io_in_wt_data_14(u_active_io_in_wt_data_14),
    .io_in_wt_data_15(u_active_io_in_wt_data_15),
    .io_in_wt_data_16(u_active_io_in_wt_data_16),
    .io_in_wt_data_17(u_active_io_in_wt_data_17),
    .io_in_wt_data_18(u_active_io_in_wt_data_18),
    .io_in_wt_data_19(u_active_io_in_wt_data_19),
    .io_in_wt_data_20(u_active_io_in_wt_data_20),
    .io_in_wt_data_21(u_active_io_in_wt_data_21),
    .io_in_wt_data_22(u_active_io_in_wt_data_22),
    .io_in_wt_data_23(u_active_io_in_wt_data_23),
    .io_in_wt_data_24(u_active_io_in_wt_data_24),
    .io_in_wt_data_25(u_active_io_in_wt_data_25),
    .io_in_wt_data_26(u_active_io_in_wt_data_26),
    .io_in_wt_data_27(u_active_io_in_wt_data_27),
    .io_in_wt_data_28(u_active_io_in_wt_data_28),
    .io_in_wt_data_29(u_active_io_in_wt_data_29),
    .io_in_wt_data_30(u_active_io_in_wt_data_30),
    .io_in_wt_data_31(u_active_io_in_wt_data_31),
    .io_in_wt_data_32(u_active_io_in_wt_data_32),
    .io_in_wt_data_33(u_active_io_in_wt_data_33),
    .io_in_wt_data_34(u_active_io_in_wt_data_34),
    .io_in_wt_data_35(u_active_io_in_wt_data_35),
    .io_in_wt_data_36(u_active_io_in_wt_data_36),
    .io_in_wt_data_37(u_active_io_in_wt_data_37),
    .io_in_wt_data_38(u_active_io_in_wt_data_38),
    .io_in_wt_data_39(u_active_io_in_wt_data_39),
    .io_in_wt_data_40(u_active_io_in_wt_data_40),
    .io_in_wt_data_41(u_active_io_in_wt_data_41),
    .io_in_wt_data_42(u_active_io_in_wt_data_42),
    .io_in_wt_data_43(u_active_io_in_wt_data_43),
    .io_in_wt_data_44(u_active_io_in_wt_data_44),
    .io_in_wt_data_45(u_active_io_in_wt_data_45),
    .io_in_wt_data_46(u_active_io_in_wt_data_46),
    .io_in_wt_data_47(u_active_io_in_wt_data_47),
    .io_in_wt_data_48(u_active_io_in_wt_data_48),
    .io_in_wt_data_49(u_active_io_in_wt_data_49),
    .io_in_wt_data_50(u_active_io_in_wt_data_50),
    .io_in_wt_data_51(u_active_io_in_wt_data_51),
    .io_in_wt_data_52(u_active_io_in_wt_data_52),
    .io_in_wt_data_53(u_active_io_in_wt_data_53),
    .io_in_wt_data_54(u_active_io_in_wt_data_54),
    .io_in_wt_data_55(u_active_io_in_wt_data_55),
    .io_in_wt_data_56(u_active_io_in_wt_data_56),
    .io_in_wt_data_57(u_active_io_in_wt_data_57),
    .io_in_wt_data_58(u_active_io_in_wt_data_58),
    .io_in_wt_data_59(u_active_io_in_wt_data_59),
    .io_in_wt_data_60(u_active_io_in_wt_data_60),
    .io_in_wt_data_61(u_active_io_in_wt_data_61),
    .io_in_wt_data_62(u_active_io_in_wt_data_62),
    .io_in_wt_data_63(u_active_io_in_wt_data_63),
    .io_in_wt_data_64(u_active_io_in_wt_data_64),
    .io_in_wt_data_65(u_active_io_in_wt_data_65),
    .io_in_wt_data_66(u_active_io_in_wt_data_66),
    .io_in_wt_data_67(u_active_io_in_wt_data_67),
    .io_in_wt_data_68(u_active_io_in_wt_data_68),
    .io_in_wt_data_69(u_active_io_in_wt_data_69),
    .io_in_wt_data_70(u_active_io_in_wt_data_70),
    .io_in_wt_data_71(u_active_io_in_wt_data_71),
    .io_in_wt_data_72(u_active_io_in_wt_data_72),
    .io_in_wt_data_73(u_active_io_in_wt_data_73),
    .io_in_wt_data_74(u_active_io_in_wt_data_74),
    .io_in_wt_data_75(u_active_io_in_wt_data_75),
    .io_in_wt_data_76(u_active_io_in_wt_data_76),
    .io_in_wt_data_77(u_active_io_in_wt_data_77),
    .io_in_wt_data_78(u_active_io_in_wt_data_78),
    .io_in_wt_data_79(u_active_io_in_wt_data_79),
    .io_in_wt_data_80(u_active_io_in_wt_data_80),
    .io_in_wt_data_81(u_active_io_in_wt_data_81),
    .io_in_wt_data_82(u_active_io_in_wt_data_82),
    .io_in_wt_data_83(u_active_io_in_wt_data_83),
    .io_in_wt_data_84(u_active_io_in_wt_data_84),
    .io_in_wt_data_85(u_active_io_in_wt_data_85),
    .io_in_wt_data_86(u_active_io_in_wt_data_86),
    .io_in_wt_data_87(u_active_io_in_wt_data_87),
    .io_in_wt_data_88(u_active_io_in_wt_data_88),
    .io_in_wt_data_89(u_active_io_in_wt_data_89),
    .io_in_wt_data_90(u_active_io_in_wt_data_90),
    .io_in_wt_data_91(u_active_io_in_wt_data_91),
    .io_in_wt_data_92(u_active_io_in_wt_data_92),
    .io_in_wt_data_93(u_active_io_in_wt_data_93),
    .io_in_wt_data_94(u_active_io_in_wt_data_94),
    .io_in_wt_data_95(u_active_io_in_wt_data_95),
    .io_in_wt_data_96(u_active_io_in_wt_data_96),
    .io_in_wt_data_97(u_active_io_in_wt_data_97),
    .io_in_wt_data_98(u_active_io_in_wt_data_98),
    .io_in_wt_data_99(u_active_io_in_wt_data_99),
    .io_in_wt_data_100(u_active_io_in_wt_data_100),
    .io_in_wt_data_101(u_active_io_in_wt_data_101),
    .io_in_wt_data_102(u_active_io_in_wt_data_102),
    .io_in_wt_data_103(u_active_io_in_wt_data_103),
    .io_in_wt_data_104(u_active_io_in_wt_data_104),
    .io_in_wt_data_105(u_active_io_in_wt_data_105),
    .io_in_wt_data_106(u_active_io_in_wt_data_106),
    .io_in_wt_data_107(u_active_io_in_wt_data_107),
    .io_in_wt_data_108(u_active_io_in_wt_data_108),
    .io_in_wt_data_109(u_active_io_in_wt_data_109),
    .io_in_wt_data_110(u_active_io_in_wt_data_110),
    .io_in_wt_data_111(u_active_io_in_wt_data_111),
    .io_in_wt_data_112(u_active_io_in_wt_data_112),
    .io_in_wt_data_113(u_active_io_in_wt_data_113),
    .io_in_wt_data_114(u_active_io_in_wt_data_114),
    .io_in_wt_data_115(u_active_io_in_wt_data_115),
    .io_in_wt_data_116(u_active_io_in_wt_data_116),
    .io_in_wt_data_117(u_active_io_in_wt_data_117),
    .io_in_wt_data_118(u_active_io_in_wt_data_118),
    .io_in_wt_data_119(u_active_io_in_wt_data_119),
    .io_in_wt_data_120(u_active_io_in_wt_data_120),
    .io_in_wt_data_121(u_active_io_in_wt_data_121),
    .io_in_wt_data_122(u_active_io_in_wt_data_122),
    .io_in_wt_data_123(u_active_io_in_wt_data_123),
    .io_in_wt_data_124(u_active_io_in_wt_data_124),
    .io_in_wt_data_125(u_active_io_in_wt_data_125),
    .io_in_wt_data_126(u_active_io_in_wt_data_126),
    .io_in_wt_data_127(u_active_io_in_wt_data_127),
    .io_in_wt_mask_0(u_active_io_in_wt_mask_0),
    .io_in_wt_mask_1(u_active_io_in_wt_mask_1),
    .io_in_wt_mask_2(u_active_io_in_wt_mask_2),
    .io_in_wt_mask_3(u_active_io_in_wt_mask_3),
    .io_in_wt_mask_4(u_active_io_in_wt_mask_4),
    .io_in_wt_mask_5(u_active_io_in_wt_mask_5),
    .io_in_wt_mask_6(u_active_io_in_wt_mask_6),
    .io_in_wt_mask_7(u_active_io_in_wt_mask_7),
    .io_in_wt_mask_8(u_active_io_in_wt_mask_8),
    .io_in_wt_mask_9(u_active_io_in_wt_mask_9),
    .io_in_wt_mask_10(u_active_io_in_wt_mask_10),
    .io_in_wt_mask_11(u_active_io_in_wt_mask_11),
    .io_in_wt_mask_12(u_active_io_in_wt_mask_12),
    .io_in_wt_mask_13(u_active_io_in_wt_mask_13),
    .io_in_wt_mask_14(u_active_io_in_wt_mask_14),
    .io_in_wt_mask_15(u_active_io_in_wt_mask_15),
    .io_in_wt_mask_16(u_active_io_in_wt_mask_16),
    .io_in_wt_mask_17(u_active_io_in_wt_mask_17),
    .io_in_wt_mask_18(u_active_io_in_wt_mask_18),
    .io_in_wt_mask_19(u_active_io_in_wt_mask_19),
    .io_in_wt_mask_20(u_active_io_in_wt_mask_20),
    .io_in_wt_mask_21(u_active_io_in_wt_mask_21),
    .io_in_wt_mask_22(u_active_io_in_wt_mask_22),
    .io_in_wt_mask_23(u_active_io_in_wt_mask_23),
    .io_in_wt_mask_24(u_active_io_in_wt_mask_24),
    .io_in_wt_mask_25(u_active_io_in_wt_mask_25),
    .io_in_wt_mask_26(u_active_io_in_wt_mask_26),
    .io_in_wt_mask_27(u_active_io_in_wt_mask_27),
    .io_in_wt_mask_28(u_active_io_in_wt_mask_28),
    .io_in_wt_mask_29(u_active_io_in_wt_mask_29),
    .io_in_wt_mask_30(u_active_io_in_wt_mask_30),
    .io_in_wt_mask_31(u_active_io_in_wt_mask_31),
    .io_in_wt_mask_32(u_active_io_in_wt_mask_32),
    .io_in_wt_mask_33(u_active_io_in_wt_mask_33),
    .io_in_wt_mask_34(u_active_io_in_wt_mask_34),
    .io_in_wt_mask_35(u_active_io_in_wt_mask_35),
    .io_in_wt_mask_36(u_active_io_in_wt_mask_36),
    .io_in_wt_mask_37(u_active_io_in_wt_mask_37),
    .io_in_wt_mask_38(u_active_io_in_wt_mask_38),
    .io_in_wt_mask_39(u_active_io_in_wt_mask_39),
    .io_in_wt_mask_40(u_active_io_in_wt_mask_40),
    .io_in_wt_mask_41(u_active_io_in_wt_mask_41),
    .io_in_wt_mask_42(u_active_io_in_wt_mask_42),
    .io_in_wt_mask_43(u_active_io_in_wt_mask_43),
    .io_in_wt_mask_44(u_active_io_in_wt_mask_44),
    .io_in_wt_mask_45(u_active_io_in_wt_mask_45),
    .io_in_wt_mask_46(u_active_io_in_wt_mask_46),
    .io_in_wt_mask_47(u_active_io_in_wt_mask_47),
    .io_in_wt_mask_48(u_active_io_in_wt_mask_48),
    .io_in_wt_mask_49(u_active_io_in_wt_mask_49),
    .io_in_wt_mask_50(u_active_io_in_wt_mask_50),
    .io_in_wt_mask_51(u_active_io_in_wt_mask_51),
    .io_in_wt_mask_52(u_active_io_in_wt_mask_52),
    .io_in_wt_mask_53(u_active_io_in_wt_mask_53),
    .io_in_wt_mask_54(u_active_io_in_wt_mask_54),
    .io_in_wt_mask_55(u_active_io_in_wt_mask_55),
    .io_in_wt_mask_56(u_active_io_in_wt_mask_56),
    .io_in_wt_mask_57(u_active_io_in_wt_mask_57),
    .io_in_wt_mask_58(u_active_io_in_wt_mask_58),
    .io_in_wt_mask_59(u_active_io_in_wt_mask_59),
    .io_in_wt_mask_60(u_active_io_in_wt_mask_60),
    .io_in_wt_mask_61(u_active_io_in_wt_mask_61),
    .io_in_wt_mask_62(u_active_io_in_wt_mask_62),
    .io_in_wt_mask_63(u_active_io_in_wt_mask_63),
    .io_in_wt_mask_64(u_active_io_in_wt_mask_64),
    .io_in_wt_mask_65(u_active_io_in_wt_mask_65),
    .io_in_wt_mask_66(u_active_io_in_wt_mask_66),
    .io_in_wt_mask_67(u_active_io_in_wt_mask_67),
    .io_in_wt_mask_68(u_active_io_in_wt_mask_68),
    .io_in_wt_mask_69(u_active_io_in_wt_mask_69),
    .io_in_wt_mask_70(u_active_io_in_wt_mask_70),
    .io_in_wt_mask_71(u_active_io_in_wt_mask_71),
    .io_in_wt_mask_72(u_active_io_in_wt_mask_72),
    .io_in_wt_mask_73(u_active_io_in_wt_mask_73),
    .io_in_wt_mask_74(u_active_io_in_wt_mask_74),
    .io_in_wt_mask_75(u_active_io_in_wt_mask_75),
    .io_in_wt_mask_76(u_active_io_in_wt_mask_76),
    .io_in_wt_mask_77(u_active_io_in_wt_mask_77),
    .io_in_wt_mask_78(u_active_io_in_wt_mask_78),
    .io_in_wt_mask_79(u_active_io_in_wt_mask_79),
    .io_in_wt_mask_80(u_active_io_in_wt_mask_80),
    .io_in_wt_mask_81(u_active_io_in_wt_mask_81),
    .io_in_wt_mask_82(u_active_io_in_wt_mask_82),
    .io_in_wt_mask_83(u_active_io_in_wt_mask_83),
    .io_in_wt_mask_84(u_active_io_in_wt_mask_84),
    .io_in_wt_mask_85(u_active_io_in_wt_mask_85),
    .io_in_wt_mask_86(u_active_io_in_wt_mask_86),
    .io_in_wt_mask_87(u_active_io_in_wt_mask_87),
    .io_in_wt_mask_88(u_active_io_in_wt_mask_88),
    .io_in_wt_mask_89(u_active_io_in_wt_mask_89),
    .io_in_wt_mask_90(u_active_io_in_wt_mask_90),
    .io_in_wt_mask_91(u_active_io_in_wt_mask_91),
    .io_in_wt_mask_92(u_active_io_in_wt_mask_92),
    .io_in_wt_mask_93(u_active_io_in_wt_mask_93),
    .io_in_wt_mask_94(u_active_io_in_wt_mask_94),
    .io_in_wt_mask_95(u_active_io_in_wt_mask_95),
    .io_in_wt_mask_96(u_active_io_in_wt_mask_96),
    .io_in_wt_mask_97(u_active_io_in_wt_mask_97),
    .io_in_wt_mask_98(u_active_io_in_wt_mask_98),
    .io_in_wt_mask_99(u_active_io_in_wt_mask_99),
    .io_in_wt_mask_100(u_active_io_in_wt_mask_100),
    .io_in_wt_mask_101(u_active_io_in_wt_mask_101),
    .io_in_wt_mask_102(u_active_io_in_wt_mask_102),
    .io_in_wt_mask_103(u_active_io_in_wt_mask_103),
    .io_in_wt_mask_104(u_active_io_in_wt_mask_104),
    .io_in_wt_mask_105(u_active_io_in_wt_mask_105),
    .io_in_wt_mask_106(u_active_io_in_wt_mask_106),
    .io_in_wt_mask_107(u_active_io_in_wt_mask_107),
    .io_in_wt_mask_108(u_active_io_in_wt_mask_108),
    .io_in_wt_mask_109(u_active_io_in_wt_mask_109),
    .io_in_wt_mask_110(u_active_io_in_wt_mask_110),
    .io_in_wt_mask_111(u_active_io_in_wt_mask_111),
    .io_in_wt_mask_112(u_active_io_in_wt_mask_112),
    .io_in_wt_mask_113(u_active_io_in_wt_mask_113),
    .io_in_wt_mask_114(u_active_io_in_wt_mask_114),
    .io_in_wt_mask_115(u_active_io_in_wt_mask_115),
    .io_in_wt_mask_116(u_active_io_in_wt_mask_116),
    .io_in_wt_mask_117(u_active_io_in_wt_mask_117),
    .io_in_wt_mask_118(u_active_io_in_wt_mask_118),
    .io_in_wt_mask_119(u_active_io_in_wt_mask_119),
    .io_in_wt_mask_120(u_active_io_in_wt_mask_120),
    .io_in_wt_mask_121(u_active_io_in_wt_mask_121),
    .io_in_wt_mask_122(u_active_io_in_wt_mask_122),
    .io_in_wt_mask_123(u_active_io_in_wt_mask_123),
    .io_in_wt_mask_124(u_active_io_in_wt_mask_124),
    .io_in_wt_mask_125(u_active_io_in_wt_mask_125),
    .io_in_wt_mask_126(u_active_io_in_wt_mask_126),
    .io_in_wt_mask_127(u_active_io_in_wt_mask_127),
    .io_in_wt_pvld(u_active_io_in_wt_pvld),
    .io_in_wt_sel_0(u_active_io_in_wt_sel_0),
    .io_dat_actv_data_0_0(u_active_io_dat_actv_data_0_0),
    .io_dat_actv_data_0_1(u_active_io_dat_actv_data_0_1),
    .io_dat_actv_data_0_2(u_active_io_dat_actv_data_0_2),
    .io_dat_actv_data_0_3(u_active_io_dat_actv_data_0_3),
    .io_dat_actv_data_0_4(u_active_io_dat_actv_data_0_4),
    .io_dat_actv_data_0_5(u_active_io_dat_actv_data_0_5),
    .io_dat_actv_data_0_6(u_active_io_dat_actv_data_0_6),
    .io_dat_actv_data_0_7(u_active_io_dat_actv_data_0_7),
    .io_dat_actv_data_0_8(u_active_io_dat_actv_data_0_8),
    .io_dat_actv_data_0_9(u_active_io_dat_actv_data_0_9),
    .io_dat_actv_data_0_10(u_active_io_dat_actv_data_0_10),
    .io_dat_actv_data_0_11(u_active_io_dat_actv_data_0_11),
    .io_dat_actv_data_0_12(u_active_io_dat_actv_data_0_12),
    .io_dat_actv_data_0_13(u_active_io_dat_actv_data_0_13),
    .io_dat_actv_data_0_14(u_active_io_dat_actv_data_0_14),
    .io_dat_actv_data_0_15(u_active_io_dat_actv_data_0_15),
    .io_dat_actv_data_0_16(u_active_io_dat_actv_data_0_16),
    .io_dat_actv_data_0_17(u_active_io_dat_actv_data_0_17),
    .io_dat_actv_data_0_18(u_active_io_dat_actv_data_0_18),
    .io_dat_actv_data_0_19(u_active_io_dat_actv_data_0_19),
    .io_dat_actv_data_0_20(u_active_io_dat_actv_data_0_20),
    .io_dat_actv_data_0_21(u_active_io_dat_actv_data_0_21),
    .io_dat_actv_data_0_22(u_active_io_dat_actv_data_0_22),
    .io_dat_actv_data_0_23(u_active_io_dat_actv_data_0_23),
    .io_dat_actv_data_0_24(u_active_io_dat_actv_data_0_24),
    .io_dat_actv_data_0_25(u_active_io_dat_actv_data_0_25),
    .io_dat_actv_data_0_26(u_active_io_dat_actv_data_0_26),
    .io_dat_actv_data_0_27(u_active_io_dat_actv_data_0_27),
    .io_dat_actv_data_0_28(u_active_io_dat_actv_data_0_28),
    .io_dat_actv_data_0_29(u_active_io_dat_actv_data_0_29),
    .io_dat_actv_data_0_30(u_active_io_dat_actv_data_0_30),
    .io_dat_actv_data_0_31(u_active_io_dat_actv_data_0_31),
    .io_dat_actv_data_0_32(u_active_io_dat_actv_data_0_32),
    .io_dat_actv_data_0_33(u_active_io_dat_actv_data_0_33),
    .io_dat_actv_data_0_34(u_active_io_dat_actv_data_0_34),
    .io_dat_actv_data_0_35(u_active_io_dat_actv_data_0_35),
    .io_dat_actv_data_0_36(u_active_io_dat_actv_data_0_36),
    .io_dat_actv_data_0_37(u_active_io_dat_actv_data_0_37),
    .io_dat_actv_data_0_38(u_active_io_dat_actv_data_0_38),
    .io_dat_actv_data_0_39(u_active_io_dat_actv_data_0_39),
    .io_dat_actv_data_0_40(u_active_io_dat_actv_data_0_40),
    .io_dat_actv_data_0_41(u_active_io_dat_actv_data_0_41),
    .io_dat_actv_data_0_42(u_active_io_dat_actv_data_0_42),
    .io_dat_actv_data_0_43(u_active_io_dat_actv_data_0_43),
    .io_dat_actv_data_0_44(u_active_io_dat_actv_data_0_44),
    .io_dat_actv_data_0_45(u_active_io_dat_actv_data_0_45),
    .io_dat_actv_data_0_46(u_active_io_dat_actv_data_0_46),
    .io_dat_actv_data_0_47(u_active_io_dat_actv_data_0_47),
    .io_dat_actv_data_0_48(u_active_io_dat_actv_data_0_48),
    .io_dat_actv_data_0_49(u_active_io_dat_actv_data_0_49),
    .io_dat_actv_data_0_50(u_active_io_dat_actv_data_0_50),
    .io_dat_actv_data_0_51(u_active_io_dat_actv_data_0_51),
    .io_dat_actv_data_0_52(u_active_io_dat_actv_data_0_52),
    .io_dat_actv_data_0_53(u_active_io_dat_actv_data_0_53),
    .io_dat_actv_data_0_54(u_active_io_dat_actv_data_0_54),
    .io_dat_actv_data_0_55(u_active_io_dat_actv_data_0_55),
    .io_dat_actv_data_0_56(u_active_io_dat_actv_data_0_56),
    .io_dat_actv_data_0_57(u_active_io_dat_actv_data_0_57),
    .io_dat_actv_data_0_58(u_active_io_dat_actv_data_0_58),
    .io_dat_actv_data_0_59(u_active_io_dat_actv_data_0_59),
    .io_dat_actv_data_0_60(u_active_io_dat_actv_data_0_60),
    .io_dat_actv_data_0_61(u_active_io_dat_actv_data_0_61),
    .io_dat_actv_data_0_62(u_active_io_dat_actv_data_0_62),
    .io_dat_actv_data_0_63(u_active_io_dat_actv_data_0_63),
    .io_dat_actv_data_0_64(u_active_io_dat_actv_data_0_64),
    .io_dat_actv_data_0_65(u_active_io_dat_actv_data_0_65),
    .io_dat_actv_data_0_66(u_active_io_dat_actv_data_0_66),
    .io_dat_actv_data_0_67(u_active_io_dat_actv_data_0_67),
    .io_dat_actv_data_0_68(u_active_io_dat_actv_data_0_68),
    .io_dat_actv_data_0_69(u_active_io_dat_actv_data_0_69),
    .io_dat_actv_data_0_70(u_active_io_dat_actv_data_0_70),
    .io_dat_actv_data_0_71(u_active_io_dat_actv_data_0_71),
    .io_dat_actv_data_0_72(u_active_io_dat_actv_data_0_72),
    .io_dat_actv_data_0_73(u_active_io_dat_actv_data_0_73),
    .io_dat_actv_data_0_74(u_active_io_dat_actv_data_0_74),
    .io_dat_actv_data_0_75(u_active_io_dat_actv_data_0_75),
    .io_dat_actv_data_0_76(u_active_io_dat_actv_data_0_76),
    .io_dat_actv_data_0_77(u_active_io_dat_actv_data_0_77),
    .io_dat_actv_data_0_78(u_active_io_dat_actv_data_0_78),
    .io_dat_actv_data_0_79(u_active_io_dat_actv_data_0_79),
    .io_dat_actv_data_0_80(u_active_io_dat_actv_data_0_80),
    .io_dat_actv_data_0_81(u_active_io_dat_actv_data_0_81),
    .io_dat_actv_data_0_82(u_active_io_dat_actv_data_0_82),
    .io_dat_actv_data_0_83(u_active_io_dat_actv_data_0_83),
    .io_dat_actv_data_0_84(u_active_io_dat_actv_data_0_84),
    .io_dat_actv_data_0_85(u_active_io_dat_actv_data_0_85),
    .io_dat_actv_data_0_86(u_active_io_dat_actv_data_0_86),
    .io_dat_actv_data_0_87(u_active_io_dat_actv_data_0_87),
    .io_dat_actv_data_0_88(u_active_io_dat_actv_data_0_88),
    .io_dat_actv_data_0_89(u_active_io_dat_actv_data_0_89),
    .io_dat_actv_data_0_90(u_active_io_dat_actv_data_0_90),
    .io_dat_actv_data_0_91(u_active_io_dat_actv_data_0_91),
    .io_dat_actv_data_0_92(u_active_io_dat_actv_data_0_92),
    .io_dat_actv_data_0_93(u_active_io_dat_actv_data_0_93),
    .io_dat_actv_data_0_94(u_active_io_dat_actv_data_0_94),
    .io_dat_actv_data_0_95(u_active_io_dat_actv_data_0_95),
    .io_dat_actv_data_0_96(u_active_io_dat_actv_data_0_96),
    .io_dat_actv_data_0_97(u_active_io_dat_actv_data_0_97),
    .io_dat_actv_data_0_98(u_active_io_dat_actv_data_0_98),
    .io_dat_actv_data_0_99(u_active_io_dat_actv_data_0_99),
    .io_dat_actv_data_0_100(u_active_io_dat_actv_data_0_100),
    .io_dat_actv_data_0_101(u_active_io_dat_actv_data_0_101),
    .io_dat_actv_data_0_102(u_active_io_dat_actv_data_0_102),
    .io_dat_actv_data_0_103(u_active_io_dat_actv_data_0_103),
    .io_dat_actv_data_0_104(u_active_io_dat_actv_data_0_104),
    .io_dat_actv_data_0_105(u_active_io_dat_actv_data_0_105),
    .io_dat_actv_data_0_106(u_active_io_dat_actv_data_0_106),
    .io_dat_actv_data_0_107(u_active_io_dat_actv_data_0_107),
    .io_dat_actv_data_0_108(u_active_io_dat_actv_data_0_108),
    .io_dat_actv_data_0_109(u_active_io_dat_actv_data_0_109),
    .io_dat_actv_data_0_110(u_active_io_dat_actv_data_0_110),
    .io_dat_actv_data_0_111(u_active_io_dat_actv_data_0_111),
    .io_dat_actv_data_0_112(u_active_io_dat_actv_data_0_112),
    .io_dat_actv_data_0_113(u_active_io_dat_actv_data_0_113),
    .io_dat_actv_data_0_114(u_active_io_dat_actv_data_0_114),
    .io_dat_actv_data_0_115(u_active_io_dat_actv_data_0_115),
    .io_dat_actv_data_0_116(u_active_io_dat_actv_data_0_116),
    .io_dat_actv_data_0_117(u_active_io_dat_actv_data_0_117),
    .io_dat_actv_data_0_118(u_active_io_dat_actv_data_0_118),
    .io_dat_actv_data_0_119(u_active_io_dat_actv_data_0_119),
    .io_dat_actv_data_0_120(u_active_io_dat_actv_data_0_120),
    .io_dat_actv_data_0_121(u_active_io_dat_actv_data_0_121),
    .io_dat_actv_data_0_122(u_active_io_dat_actv_data_0_122),
    .io_dat_actv_data_0_123(u_active_io_dat_actv_data_0_123),
    .io_dat_actv_data_0_124(u_active_io_dat_actv_data_0_124),
    .io_dat_actv_data_0_125(u_active_io_dat_actv_data_0_125),
    .io_dat_actv_data_0_126(u_active_io_dat_actv_data_0_126),
    .io_dat_actv_data_0_127(u_active_io_dat_actv_data_0_127),
    .io_dat_actv_nz_0_0(u_active_io_dat_actv_nz_0_0),
    .io_dat_actv_nz_0_1(u_active_io_dat_actv_nz_0_1),
    .io_dat_actv_nz_0_2(u_active_io_dat_actv_nz_0_2),
    .io_dat_actv_nz_0_3(u_active_io_dat_actv_nz_0_3),
    .io_dat_actv_nz_0_4(u_active_io_dat_actv_nz_0_4),
    .io_dat_actv_nz_0_5(u_active_io_dat_actv_nz_0_5),
    .io_dat_actv_nz_0_6(u_active_io_dat_actv_nz_0_6),
    .io_dat_actv_nz_0_7(u_active_io_dat_actv_nz_0_7),
    .io_dat_actv_nz_0_8(u_active_io_dat_actv_nz_0_8),
    .io_dat_actv_nz_0_9(u_active_io_dat_actv_nz_0_9),
    .io_dat_actv_nz_0_10(u_active_io_dat_actv_nz_0_10),
    .io_dat_actv_nz_0_11(u_active_io_dat_actv_nz_0_11),
    .io_dat_actv_nz_0_12(u_active_io_dat_actv_nz_0_12),
    .io_dat_actv_nz_0_13(u_active_io_dat_actv_nz_0_13),
    .io_dat_actv_nz_0_14(u_active_io_dat_actv_nz_0_14),
    .io_dat_actv_nz_0_15(u_active_io_dat_actv_nz_0_15),
    .io_dat_actv_nz_0_16(u_active_io_dat_actv_nz_0_16),
    .io_dat_actv_nz_0_17(u_active_io_dat_actv_nz_0_17),
    .io_dat_actv_nz_0_18(u_active_io_dat_actv_nz_0_18),
    .io_dat_actv_nz_0_19(u_active_io_dat_actv_nz_0_19),
    .io_dat_actv_nz_0_20(u_active_io_dat_actv_nz_0_20),
    .io_dat_actv_nz_0_21(u_active_io_dat_actv_nz_0_21),
    .io_dat_actv_nz_0_22(u_active_io_dat_actv_nz_0_22),
    .io_dat_actv_nz_0_23(u_active_io_dat_actv_nz_0_23),
    .io_dat_actv_nz_0_24(u_active_io_dat_actv_nz_0_24),
    .io_dat_actv_nz_0_25(u_active_io_dat_actv_nz_0_25),
    .io_dat_actv_nz_0_26(u_active_io_dat_actv_nz_0_26),
    .io_dat_actv_nz_0_27(u_active_io_dat_actv_nz_0_27),
    .io_dat_actv_nz_0_28(u_active_io_dat_actv_nz_0_28),
    .io_dat_actv_nz_0_29(u_active_io_dat_actv_nz_0_29),
    .io_dat_actv_nz_0_30(u_active_io_dat_actv_nz_0_30),
    .io_dat_actv_nz_0_31(u_active_io_dat_actv_nz_0_31),
    .io_dat_actv_nz_0_32(u_active_io_dat_actv_nz_0_32),
    .io_dat_actv_nz_0_33(u_active_io_dat_actv_nz_0_33),
    .io_dat_actv_nz_0_34(u_active_io_dat_actv_nz_0_34),
    .io_dat_actv_nz_0_35(u_active_io_dat_actv_nz_0_35),
    .io_dat_actv_nz_0_36(u_active_io_dat_actv_nz_0_36),
    .io_dat_actv_nz_0_37(u_active_io_dat_actv_nz_0_37),
    .io_dat_actv_nz_0_38(u_active_io_dat_actv_nz_0_38),
    .io_dat_actv_nz_0_39(u_active_io_dat_actv_nz_0_39),
    .io_dat_actv_nz_0_40(u_active_io_dat_actv_nz_0_40),
    .io_dat_actv_nz_0_41(u_active_io_dat_actv_nz_0_41),
    .io_dat_actv_nz_0_42(u_active_io_dat_actv_nz_0_42),
    .io_dat_actv_nz_0_43(u_active_io_dat_actv_nz_0_43),
    .io_dat_actv_nz_0_44(u_active_io_dat_actv_nz_0_44),
    .io_dat_actv_nz_0_45(u_active_io_dat_actv_nz_0_45),
    .io_dat_actv_nz_0_46(u_active_io_dat_actv_nz_0_46),
    .io_dat_actv_nz_0_47(u_active_io_dat_actv_nz_0_47),
    .io_dat_actv_nz_0_48(u_active_io_dat_actv_nz_0_48),
    .io_dat_actv_nz_0_49(u_active_io_dat_actv_nz_0_49),
    .io_dat_actv_nz_0_50(u_active_io_dat_actv_nz_0_50),
    .io_dat_actv_nz_0_51(u_active_io_dat_actv_nz_0_51),
    .io_dat_actv_nz_0_52(u_active_io_dat_actv_nz_0_52),
    .io_dat_actv_nz_0_53(u_active_io_dat_actv_nz_0_53),
    .io_dat_actv_nz_0_54(u_active_io_dat_actv_nz_0_54),
    .io_dat_actv_nz_0_55(u_active_io_dat_actv_nz_0_55),
    .io_dat_actv_nz_0_56(u_active_io_dat_actv_nz_0_56),
    .io_dat_actv_nz_0_57(u_active_io_dat_actv_nz_0_57),
    .io_dat_actv_nz_0_58(u_active_io_dat_actv_nz_0_58),
    .io_dat_actv_nz_0_59(u_active_io_dat_actv_nz_0_59),
    .io_dat_actv_nz_0_60(u_active_io_dat_actv_nz_0_60),
    .io_dat_actv_nz_0_61(u_active_io_dat_actv_nz_0_61),
    .io_dat_actv_nz_0_62(u_active_io_dat_actv_nz_0_62),
    .io_dat_actv_nz_0_63(u_active_io_dat_actv_nz_0_63),
    .io_dat_actv_nz_0_64(u_active_io_dat_actv_nz_0_64),
    .io_dat_actv_nz_0_65(u_active_io_dat_actv_nz_0_65),
    .io_dat_actv_nz_0_66(u_active_io_dat_actv_nz_0_66),
    .io_dat_actv_nz_0_67(u_active_io_dat_actv_nz_0_67),
    .io_dat_actv_nz_0_68(u_active_io_dat_actv_nz_0_68),
    .io_dat_actv_nz_0_69(u_active_io_dat_actv_nz_0_69),
    .io_dat_actv_nz_0_70(u_active_io_dat_actv_nz_0_70),
    .io_dat_actv_nz_0_71(u_active_io_dat_actv_nz_0_71),
    .io_dat_actv_nz_0_72(u_active_io_dat_actv_nz_0_72),
    .io_dat_actv_nz_0_73(u_active_io_dat_actv_nz_0_73),
    .io_dat_actv_nz_0_74(u_active_io_dat_actv_nz_0_74),
    .io_dat_actv_nz_0_75(u_active_io_dat_actv_nz_0_75),
    .io_dat_actv_nz_0_76(u_active_io_dat_actv_nz_0_76),
    .io_dat_actv_nz_0_77(u_active_io_dat_actv_nz_0_77),
    .io_dat_actv_nz_0_78(u_active_io_dat_actv_nz_0_78),
    .io_dat_actv_nz_0_79(u_active_io_dat_actv_nz_0_79),
    .io_dat_actv_nz_0_80(u_active_io_dat_actv_nz_0_80),
    .io_dat_actv_nz_0_81(u_active_io_dat_actv_nz_0_81),
    .io_dat_actv_nz_0_82(u_active_io_dat_actv_nz_0_82),
    .io_dat_actv_nz_0_83(u_active_io_dat_actv_nz_0_83),
    .io_dat_actv_nz_0_84(u_active_io_dat_actv_nz_0_84),
    .io_dat_actv_nz_0_85(u_active_io_dat_actv_nz_0_85),
    .io_dat_actv_nz_0_86(u_active_io_dat_actv_nz_0_86),
    .io_dat_actv_nz_0_87(u_active_io_dat_actv_nz_0_87),
    .io_dat_actv_nz_0_88(u_active_io_dat_actv_nz_0_88),
    .io_dat_actv_nz_0_89(u_active_io_dat_actv_nz_0_89),
    .io_dat_actv_nz_0_90(u_active_io_dat_actv_nz_0_90),
    .io_dat_actv_nz_0_91(u_active_io_dat_actv_nz_0_91),
    .io_dat_actv_nz_0_92(u_active_io_dat_actv_nz_0_92),
    .io_dat_actv_nz_0_93(u_active_io_dat_actv_nz_0_93),
    .io_dat_actv_nz_0_94(u_active_io_dat_actv_nz_0_94),
    .io_dat_actv_nz_0_95(u_active_io_dat_actv_nz_0_95),
    .io_dat_actv_nz_0_96(u_active_io_dat_actv_nz_0_96),
    .io_dat_actv_nz_0_97(u_active_io_dat_actv_nz_0_97),
    .io_dat_actv_nz_0_98(u_active_io_dat_actv_nz_0_98),
    .io_dat_actv_nz_0_99(u_active_io_dat_actv_nz_0_99),
    .io_dat_actv_nz_0_100(u_active_io_dat_actv_nz_0_100),
    .io_dat_actv_nz_0_101(u_active_io_dat_actv_nz_0_101),
    .io_dat_actv_nz_0_102(u_active_io_dat_actv_nz_0_102),
    .io_dat_actv_nz_0_103(u_active_io_dat_actv_nz_0_103),
    .io_dat_actv_nz_0_104(u_active_io_dat_actv_nz_0_104),
    .io_dat_actv_nz_0_105(u_active_io_dat_actv_nz_0_105),
    .io_dat_actv_nz_0_106(u_active_io_dat_actv_nz_0_106),
    .io_dat_actv_nz_0_107(u_active_io_dat_actv_nz_0_107),
    .io_dat_actv_nz_0_108(u_active_io_dat_actv_nz_0_108),
    .io_dat_actv_nz_0_109(u_active_io_dat_actv_nz_0_109),
    .io_dat_actv_nz_0_110(u_active_io_dat_actv_nz_0_110),
    .io_dat_actv_nz_0_111(u_active_io_dat_actv_nz_0_111),
    .io_dat_actv_nz_0_112(u_active_io_dat_actv_nz_0_112),
    .io_dat_actv_nz_0_113(u_active_io_dat_actv_nz_0_113),
    .io_dat_actv_nz_0_114(u_active_io_dat_actv_nz_0_114),
    .io_dat_actv_nz_0_115(u_active_io_dat_actv_nz_0_115),
    .io_dat_actv_nz_0_116(u_active_io_dat_actv_nz_0_116),
    .io_dat_actv_nz_0_117(u_active_io_dat_actv_nz_0_117),
    .io_dat_actv_nz_0_118(u_active_io_dat_actv_nz_0_118),
    .io_dat_actv_nz_0_119(u_active_io_dat_actv_nz_0_119),
    .io_dat_actv_nz_0_120(u_active_io_dat_actv_nz_0_120),
    .io_dat_actv_nz_0_121(u_active_io_dat_actv_nz_0_121),
    .io_dat_actv_nz_0_122(u_active_io_dat_actv_nz_0_122),
    .io_dat_actv_nz_0_123(u_active_io_dat_actv_nz_0_123),
    .io_dat_actv_nz_0_124(u_active_io_dat_actv_nz_0_124),
    .io_dat_actv_nz_0_125(u_active_io_dat_actv_nz_0_125),
    .io_dat_actv_nz_0_126(u_active_io_dat_actv_nz_0_126),
    .io_dat_actv_nz_0_127(u_active_io_dat_actv_nz_0_127),
    .io_dat_actv_pvld_0_0(u_active_io_dat_actv_pvld_0_0),
    .io_dat_actv_pvld_0_1(u_active_io_dat_actv_pvld_0_1),
    .io_dat_actv_pvld_0_2(u_active_io_dat_actv_pvld_0_2),
    .io_dat_actv_pvld_0_3(u_active_io_dat_actv_pvld_0_3),
    .io_dat_actv_pvld_0_4(u_active_io_dat_actv_pvld_0_4),
    .io_dat_actv_pvld_0_5(u_active_io_dat_actv_pvld_0_5),
    .io_dat_actv_pvld_0_6(u_active_io_dat_actv_pvld_0_6),
    .io_dat_actv_pvld_0_7(u_active_io_dat_actv_pvld_0_7),
    .io_dat_actv_pvld_0_8(u_active_io_dat_actv_pvld_0_8),
    .io_dat_actv_pvld_0_9(u_active_io_dat_actv_pvld_0_9),
    .io_dat_actv_pvld_0_10(u_active_io_dat_actv_pvld_0_10),
    .io_dat_actv_pvld_0_11(u_active_io_dat_actv_pvld_0_11),
    .io_dat_actv_pvld_0_12(u_active_io_dat_actv_pvld_0_12),
    .io_dat_actv_pvld_0_13(u_active_io_dat_actv_pvld_0_13),
    .io_dat_actv_pvld_0_14(u_active_io_dat_actv_pvld_0_14),
    .io_dat_actv_pvld_0_15(u_active_io_dat_actv_pvld_0_15),
    .io_dat_actv_pvld_0_16(u_active_io_dat_actv_pvld_0_16),
    .io_dat_actv_pvld_0_17(u_active_io_dat_actv_pvld_0_17),
    .io_dat_actv_pvld_0_18(u_active_io_dat_actv_pvld_0_18),
    .io_dat_actv_pvld_0_19(u_active_io_dat_actv_pvld_0_19),
    .io_dat_actv_pvld_0_20(u_active_io_dat_actv_pvld_0_20),
    .io_dat_actv_pvld_0_21(u_active_io_dat_actv_pvld_0_21),
    .io_dat_actv_pvld_0_22(u_active_io_dat_actv_pvld_0_22),
    .io_dat_actv_pvld_0_23(u_active_io_dat_actv_pvld_0_23),
    .io_dat_actv_pvld_0_24(u_active_io_dat_actv_pvld_0_24),
    .io_dat_actv_pvld_0_25(u_active_io_dat_actv_pvld_0_25),
    .io_dat_actv_pvld_0_26(u_active_io_dat_actv_pvld_0_26),
    .io_dat_actv_pvld_0_27(u_active_io_dat_actv_pvld_0_27),
    .io_dat_actv_pvld_0_28(u_active_io_dat_actv_pvld_0_28),
    .io_dat_actv_pvld_0_29(u_active_io_dat_actv_pvld_0_29),
    .io_dat_actv_pvld_0_30(u_active_io_dat_actv_pvld_0_30),
    .io_dat_actv_pvld_0_31(u_active_io_dat_actv_pvld_0_31),
    .io_dat_actv_pvld_0_32(u_active_io_dat_actv_pvld_0_32),
    .io_dat_actv_pvld_0_33(u_active_io_dat_actv_pvld_0_33),
    .io_dat_actv_pvld_0_34(u_active_io_dat_actv_pvld_0_34),
    .io_dat_actv_pvld_0_35(u_active_io_dat_actv_pvld_0_35),
    .io_dat_actv_pvld_0_36(u_active_io_dat_actv_pvld_0_36),
    .io_dat_actv_pvld_0_37(u_active_io_dat_actv_pvld_0_37),
    .io_dat_actv_pvld_0_38(u_active_io_dat_actv_pvld_0_38),
    .io_dat_actv_pvld_0_39(u_active_io_dat_actv_pvld_0_39),
    .io_dat_actv_pvld_0_40(u_active_io_dat_actv_pvld_0_40),
    .io_dat_actv_pvld_0_41(u_active_io_dat_actv_pvld_0_41),
    .io_dat_actv_pvld_0_42(u_active_io_dat_actv_pvld_0_42),
    .io_dat_actv_pvld_0_43(u_active_io_dat_actv_pvld_0_43),
    .io_dat_actv_pvld_0_44(u_active_io_dat_actv_pvld_0_44),
    .io_dat_actv_pvld_0_45(u_active_io_dat_actv_pvld_0_45),
    .io_dat_actv_pvld_0_46(u_active_io_dat_actv_pvld_0_46),
    .io_dat_actv_pvld_0_47(u_active_io_dat_actv_pvld_0_47),
    .io_dat_actv_pvld_0_48(u_active_io_dat_actv_pvld_0_48),
    .io_dat_actv_pvld_0_49(u_active_io_dat_actv_pvld_0_49),
    .io_dat_actv_pvld_0_50(u_active_io_dat_actv_pvld_0_50),
    .io_dat_actv_pvld_0_51(u_active_io_dat_actv_pvld_0_51),
    .io_dat_actv_pvld_0_52(u_active_io_dat_actv_pvld_0_52),
    .io_dat_actv_pvld_0_53(u_active_io_dat_actv_pvld_0_53),
    .io_dat_actv_pvld_0_54(u_active_io_dat_actv_pvld_0_54),
    .io_dat_actv_pvld_0_55(u_active_io_dat_actv_pvld_0_55),
    .io_dat_actv_pvld_0_56(u_active_io_dat_actv_pvld_0_56),
    .io_dat_actv_pvld_0_57(u_active_io_dat_actv_pvld_0_57),
    .io_dat_actv_pvld_0_58(u_active_io_dat_actv_pvld_0_58),
    .io_dat_actv_pvld_0_59(u_active_io_dat_actv_pvld_0_59),
    .io_dat_actv_pvld_0_60(u_active_io_dat_actv_pvld_0_60),
    .io_dat_actv_pvld_0_61(u_active_io_dat_actv_pvld_0_61),
    .io_dat_actv_pvld_0_62(u_active_io_dat_actv_pvld_0_62),
    .io_dat_actv_pvld_0_63(u_active_io_dat_actv_pvld_0_63),
    .io_dat_actv_pvld_0_64(u_active_io_dat_actv_pvld_0_64),
    .io_dat_actv_pvld_0_65(u_active_io_dat_actv_pvld_0_65),
    .io_dat_actv_pvld_0_66(u_active_io_dat_actv_pvld_0_66),
    .io_dat_actv_pvld_0_67(u_active_io_dat_actv_pvld_0_67),
    .io_dat_actv_pvld_0_68(u_active_io_dat_actv_pvld_0_68),
    .io_dat_actv_pvld_0_69(u_active_io_dat_actv_pvld_0_69),
    .io_dat_actv_pvld_0_70(u_active_io_dat_actv_pvld_0_70),
    .io_dat_actv_pvld_0_71(u_active_io_dat_actv_pvld_0_71),
    .io_dat_actv_pvld_0_72(u_active_io_dat_actv_pvld_0_72),
    .io_dat_actv_pvld_0_73(u_active_io_dat_actv_pvld_0_73),
    .io_dat_actv_pvld_0_74(u_active_io_dat_actv_pvld_0_74),
    .io_dat_actv_pvld_0_75(u_active_io_dat_actv_pvld_0_75),
    .io_dat_actv_pvld_0_76(u_active_io_dat_actv_pvld_0_76),
    .io_dat_actv_pvld_0_77(u_active_io_dat_actv_pvld_0_77),
    .io_dat_actv_pvld_0_78(u_active_io_dat_actv_pvld_0_78),
    .io_dat_actv_pvld_0_79(u_active_io_dat_actv_pvld_0_79),
    .io_dat_actv_pvld_0_80(u_active_io_dat_actv_pvld_0_80),
    .io_dat_actv_pvld_0_81(u_active_io_dat_actv_pvld_0_81),
    .io_dat_actv_pvld_0_82(u_active_io_dat_actv_pvld_0_82),
    .io_dat_actv_pvld_0_83(u_active_io_dat_actv_pvld_0_83),
    .io_dat_actv_pvld_0_84(u_active_io_dat_actv_pvld_0_84),
    .io_dat_actv_pvld_0_85(u_active_io_dat_actv_pvld_0_85),
    .io_dat_actv_pvld_0_86(u_active_io_dat_actv_pvld_0_86),
    .io_dat_actv_pvld_0_87(u_active_io_dat_actv_pvld_0_87),
    .io_dat_actv_pvld_0_88(u_active_io_dat_actv_pvld_0_88),
    .io_dat_actv_pvld_0_89(u_active_io_dat_actv_pvld_0_89),
    .io_dat_actv_pvld_0_90(u_active_io_dat_actv_pvld_0_90),
    .io_dat_actv_pvld_0_91(u_active_io_dat_actv_pvld_0_91),
    .io_dat_actv_pvld_0_92(u_active_io_dat_actv_pvld_0_92),
    .io_dat_actv_pvld_0_93(u_active_io_dat_actv_pvld_0_93),
    .io_dat_actv_pvld_0_94(u_active_io_dat_actv_pvld_0_94),
    .io_dat_actv_pvld_0_95(u_active_io_dat_actv_pvld_0_95),
    .io_dat_actv_pvld_0_96(u_active_io_dat_actv_pvld_0_96),
    .io_dat_actv_pvld_0_97(u_active_io_dat_actv_pvld_0_97),
    .io_dat_actv_pvld_0_98(u_active_io_dat_actv_pvld_0_98),
    .io_dat_actv_pvld_0_99(u_active_io_dat_actv_pvld_0_99),
    .io_dat_actv_pvld_0_100(u_active_io_dat_actv_pvld_0_100),
    .io_dat_actv_pvld_0_101(u_active_io_dat_actv_pvld_0_101),
    .io_dat_actv_pvld_0_102(u_active_io_dat_actv_pvld_0_102),
    .io_dat_actv_pvld_0_103(u_active_io_dat_actv_pvld_0_103),
    .io_dat_actv_pvld_0_104(u_active_io_dat_actv_pvld_0_104),
    .io_dat_actv_pvld_0_105(u_active_io_dat_actv_pvld_0_105),
    .io_dat_actv_pvld_0_106(u_active_io_dat_actv_pvld_0_106),
    .io_dat_actv_pvld_0_107(u_active_io_dat_actv_pvld_0_107),
    .io_dat_actv_pvld_0_108(u_active_io_dat_actv_pvld_0_108),
    .io_dat_actv_pvld_0_109(u_active_io_dat_actv_pvld_0_109),
    .io_dat_actv_pvld_0_110(u_active_io_dat_actv_pvld_0_110),
    .io_dat_actv_pvld_0_111(u_active_io_dat_actv_pvld_0_111),
    .io_dat_actv_pvld_0_112(u_active_io_dat_actv_pvld_0_112),
    .io_dat_actv_pvld_0_113(u_active_io_dat_actv_pvld_0_113),
    .io_dat_actv_pvld_0_114(u_active_io_dat_actv_pvld_0_114),
    .io_dat_actv_pvld_0_115(u_active_io_dat_actv_pvld_0_115),
    .io_dat_actv_pvld_0_116(u_active_io_dat_actv_pvld_0_116),
    .io_dat_actv_pvld_0_117(u_active_io_dat_actv_pvld_0_117),
    .io_dat_actv_pvld_0_118(u_active_io_dat_actv_pvld_0_118),
    .io_dat_actv_pvld_0_119(u_active_io_dat_actv_pvld_0_119),
    .io_dat_actv_pvld_0_120(u_active_io_dat_actv_pvld_0_120),
    .io_dat_actv_pvld_0_121(u_active_io_dat_actv_pvld_0_121),
    .io_dat_actv_pvld_0_122(u_active_io_dat_actv_pvld_0_122),
    .io_dat_actv_pvld_0_123(u_active_io_dat_actv_pvld_0_123),
    .io_dat_actv_pvld_0_124(u_active_io_dat_actv_pvld_0_124),
    .io_dat_actv_pvld_0_125(u_active_io_dat_actv_pvld_0_125),
    .io_dat_actv_pvld_0_126(u_active_io_dat_actv_pvld_0_126),
    .io_dat_actv_pvld_0_127(u_active_io_dat_actv_pvld_0_127),
    .io_wt_actv_data_0_0(u_active_io_wt_actv_data_0_0),
    .io_wt_actv_data_0_1(u_active_io_wt_actv_data_0_1),
    .io_wt_actv_data_0_2(u_active_io_wt_actv_data_0_2),
    .io_wt_actv_data_0_3(u_active_io_wt_actv_data_0_3),
    .io_wt_actv_data_0_4(u_active_io_wt_actv_data_0_4),
    .io_wt_actv_data_0_5(u_active_io_wt_actv_data_0_5),
    .io_wt_actv_data_0_6(u_active_io_wt_actv_data_0_6),
    .io_wt_actv_data_0_7(u_active_io_wt_actv_data_0_7),
    .io_wt_actv_data_0_8(u_active_io_wt_actv_data_0_8),
    .io_wt_actv_data_0_9(u_active_io_wt_actv_data_0_9),
    .io_wt_actv_data_0_10(u_active_io_wt_actv_data_0_10),
    .io_wt_actv_data_0_11(u_active_io_wt_actv_data_0_11),
    .io_wt_actv_data_0_12(u_active_io_wt_actv_data_0_12),
    .io_wt_actv_data_0_13(u_active_io_wt_actv_data_0_13),
    .io_wt_actv_data_0_14(u_active_io_wt_actv_data_0_14),
    .io_wt_actv_data_0_15(u_active_io_wt_actv_data_0_15),
    .io_wt_actv_data_0_16(u_active_io_wt_actv_data_0_16),
    .io_wt_actv_data_0_17(u_active_io_wt_actv_data_0_17),
    .io_wt_actv_data_0_18(u_active_io_wt_actv_data_0_18),
    .io_wt_actv_data_0_19(u_active_io_wt_actv_data_0_19),
    .io_wt_actv_data_0_20(u_active_io_wt_actv_data_0_20),
    .io_wt_actv_data_0_21(u_active_io_wt_actv_data_0_21),
    .io_wt_actv_data_0_22(u_active_io_wt_actv_data_0_22),
    .io_wt_actv_data_0_23(u_active_io_wt_actv_data_0_23),
    .io_wt_actv_data_0_24(u_active_io_wt_actv_data_0_24),
    .io_wt_actv_data_0_25(u_active_io_wt_actv_data_0_25),
    .io_wt_actv_data_0_26(u_active_io_wt_actv_data_0_26),
    .io_wt_actv_data_0_27(u_active_io_wt_actv_data_0_27),
    .io_wt_actv_data_0_28(u_active_io_wt_actv_data_0_28),
    .io_wt_actv_data_0_29(u_active_io_wt_actv_data_0_29),
    .io_wt_actv_data_0_30(u_active_io_wt_actv_data_0_30),
    .io_wt_actv_data_0_31(u_active_io_wt_actv_data_0_31),
    .io_wt_actv_data_0_32(u_active_io_wt_actv_data_0_32),
    .io_wt_actv_data_0_33(u_active_io_wt_actv_data_0_33),
    .io_wt_actv_data_0_34(u_active_io_wt_actv_data_0_34),
    .io_wt_actv_data_0_35(u_active_io_wt_actv_data_0_35),
    .io_wt_actv_data_0_36(u_active_io_wt_actv_data_0_36),
    .io_wt_actv_data_0_37(u_active_io_wt_actv_data_0_37),
    .io_wt_actv_data_0_38(u_active_io_wt_actv_data_0_38),
    .io_wt_actv_data_0_39(u_active_io_wt_actv_data_0_39),
    .io_wt_actv_data_0_40(u_active_io_wt_actv_data_0_40),
    .io_wt_actv_data_0_41(u_active_io_wt_actv_data_0_41),
    .io_wt_actv_data_0_42(u_active_io_wt_actv_data_0_42),
    .io_wt_actv_data_0_43(u_active_io_wt_actv_data_0_43),
    .io_wt_actv_data_0_44(u_active_io_wt_actv_data_0_44),
    .io_wt_actv_data_0_45(u_active_io_wt_actv_data_0_45),
    .io_wt_actv_data_0_46(u_active_io_wt_actv_data_0_46),
    .io_wt_actv_data_0_47(u_active_io_wt_actv_data_0_47),
    .io_wt_actv_data_0_48(u_active_io_wt_actv_data_0_48),
    .io_wt_actv_data_0_49(u_active_io_wt_actv_data_0_49),
    .io_wt_actv_data_0_50(u_active_io_wt_actv_data_0_50),
    .io_wt_actv_data_0_51(u_active_io_wt_actv_data_0_51),
    .io_wt_actv_data_0_52(u_active_io_wt_actv_data_0_52),
    .io_wt_actv_data_0_53(u_active_io_wt_actv_data_0_53),
    .io_wt_actv_data_0_54(u_active_io_wt_actv_data_0_54),
    .io_wt_actv_data_0_55(u_active_io_wt_actv_data_0_55),
    .io_wt_actv_data_0_56(u_active_io_wt_actv_data_0_56),
    .io_wt_actv_data_0_57(u_active_io_wt_actv_data_0_57),
    .io_wt_actv_data_0_58(u_active_io_wt_actv_data_0_58),
    .io_wt_actv_data_0_59(u_active_io_wt_actv_data_0_59),
    .io_wt_actv_data_0_60(u_active_io_wt_actv_data_0_60),
    .io_wt_actv_data_0_61(u_active_io_wt_actv_data_0_61),
    .io_wt_actv_data_0_62(u_active_io_wt_actv_data_0_62),
    .io_wt_actv_data_0_63(u_active_io_wt_actv_data_0_63),
    .io_wt_actv_data_0_64(u_active_io_wt_actv_data_0_64),
    .io_wt_actv_data_0_65(u_active_io_wt_actv_data_0_65),
    .io_wt_actv_data_0_66(u_active_io_wt_actv_data_0_66),
    .io_wt_actv_data_0_67(u_active_io_wt_actv_data_0_67),
    .io_wt_actv_data_0_68(u_active_io_wt_actv_data_0_68),
    .io_wt_actv_data_0_69(u_active_io_wt_actv_data_0_69),
    .io_wt_actv_data_0_70(u_active_io_wt_actv_data_0_70),
    .io_wt_actv_data_0_71(u_active_io_wt_actv_data_0_71),
    .io_wt_actv_data_0_72(u_active_io_wt_actv_data_0_72),
    .io_wt_actv_data_0_73(u_active_io_wt_actv_data_0_73),
    .io_wt_actv_data_0_74(u_active_io_wt_actv_data_0_74),
    .io_wt_actv_data_0_75(u_active_io_wt_actv_data_0_75),
    .io_wt_actv_data_0_76(u_active_io_wt_actv_data_0_76),
    .io_wt_actv_data_0_77(u_active_io_wt_actv_data_0_77),
    .io_wt_actv_data_0_78(u_active_io_wt_actv_data_0_78),
    .io_wt_actv_data_0_79(u_active_io_wt_actv_data_0_79),
    .io_wt_actv_data_0_80(u_active_io_wt_actv_data_0_80),
    .io_wt_actv_data_0_81(u_active_io_wt_actv_data_0_81),
    .io_wt_actv_data_0_82(u_active_io_wt_actv_data_0_82),
    .io_wt_actv_data_0_83(u_active_io_wt_actv_data_0_83),
    .io_wt_actv_data_0_84(u_active_io_wt_actv_data_0_84),
    .io_wt_actv_data_0_85(u_active_io_wt_actv_data_0_85),
    .io_wt_actv_data_0_86(u_active_io_wt_actv_data_0_86),
    .io_wt_actv_data_0_87(u_active_io_wt_actv_data_0_87),
    .io_wt_actv_data_0_88(u_active_io_wt_actv_data_0_88),
    .io_wt_actv_data_0_89(u_active_io_wt_actv_data_0_89),
    .io_wt_actv_data_0_90(u_active_io_wt_actv_data_0_90),
    .io_wt_actv_data_0_91(u_active_io_wt_actv_data_0_91),
    .io_wt_actv_data_0_92(u_active_io_wt_actv_data_0_92),
    .io_wt_actv_data_0_93(u_active_io_wt_actv_data_0_93),
    .io_wt_actv_data_0_94(u_active_io_wt_actv_data_0_94),
    .io_wt_actv_data_0_95(u_active_io_wt_actv_data_0_95),
    .io_wt_actv_data_0_96(u_active_io_wt_actv_data_0_96),
    .io_wt_actv_data_0_97(u_active_io_wt_actv_data_0_97),
    .io_wt_actv_data_0_98(u_active_io_wt_actv_data_0_98),
    .io_wt_actv_data_0_99(u_active_io_wt_actv_data_0_99),
    .io_wt_actv_data_0_100(u_active_io_wt_actv_data_0_100),
    .io_wt_actv_data_0_101(u_active_io_wt_actv_data_0_101),
    .io_wt_actv_data_0_102(u_active_io_wt_actv_data_0_102),
    .io_wt_actv_data_0_103(u_active_io_wt_actv_data_0_103),
    .io_wt_actv_data_0_104(u_active_io_wt_actv_data_0_104),
    .io_wt_actv_data_0_105(u_active_io_wt_actv_data_0_105),
    .io_wt_actv_data_0_106(u_active_io_wt_actv_data_0_106),
    .io_wt_actv_data_0_107(u_active_io_wt_actv_data_0_107),
    .io_wt_actv_data_0_108(u_active_io_wt_actv_data_0_108),
    .io_wt_actv_data_0_109(u_active_io_wt_actv_data_0_109),
    .io_wt_actv_data_0_110(u_active_io_wt_actv_data_0_110),
    .io_wt_actv_data_0_111(u_active_io_wt_actv_data_0_111),
    .io_wt_actv_data_0_112(u_active_io_wt_actv_data_0_112),
    .io_wt_actv_data_0_113(u_active_io_wt_actv_data_0_113),
    .io_wt_actv_data_0_114(u_active_io_wt_actv_data_0_114),
    .io_wt_actv_data_0_115(u_active_io_wt_actv_data_0_115),
    .io_wt_actv_data_0_116(u_active_io_wt_actv_data_0_116),
    .io_wt_actv_data_0_117(u_active_io_wt_actv_data_0_117),
    .io_wt_actv_data_0_118(u_active_io_wt_actv_data_0_118),
    .io_wt_actv_data_0_119(u_active_io_wt_actv_data_0_119),
    .io_wt_actv_data_0_120(u_active_io_wt_actv_data_0_120),
    .io_wt_actv_data_0_121(u_active_io_wt_actv_data_0_121),
    .io_wt_actv_data_0_122(u_active_io_wt_actv_data_0_122),
    .io_wt_actv_data_0_123(u_active_io_wt_actv_data_0_123),
    .io_wt_actv_data_0_124(u_active_io_wt_actv_data_0_124),
    .io_wt_actv_data_0_125(u_active_io_wt_actv_data_0_125),
    .io_wt_actv_data_0_126(u_active_io_wt_actv_data_0_126),
    .io_wt_actv_data_0_127(u_active_io_wt_actv_data_0_127),
    .io_wt_actv_nz_0_0(u_active_io_wt_actv_nz_0_0),
    .io_wt_actv_nz_0_1(u_active_io_wt_actv_nz_0_1),
    .io_wt_actv_nz_0_2(u_active_io_wt_actv_nz_0_2),
    .io_wt_actv_nz_0_3(u_active_io_wt_actv_nz_0_3),
    .io_wt_actv_nz_0_4(u_active_io_wt_actv_nz_0_4),
    .io_wt_actv_nz_0_5(u_active_io_wt_actv_nz_0_5),
    .io_wt_actv_nz_0_6(u_active_io_wt_actv_nz_0_6),
    .io_wt_actv_nz_0_7(u_active_io_wt_actv_nz_0_7),
    .io_wt_actv_nz_0_8(u_active_io_wt_actv_nz_0_8),
    .io_wt_actv_nz_0_9(u_active_io_wt_actv_nz_0_9),
    .io_wt_actv_nz_0_10(u_active_io_wt_actv_nz_0_10),
    .io_wt_actv_nz_0_11(u_active_io_wt_actv_nz_0_11),
    .io_wt_actv_nz_0_12(u_active_io_wt_actv_nz_0_12),
    .io_wt_actv_nz_0_13(u_active_io_wt_actv_nz_0_13),
    .io_wt_actv_nz_0_14(u_active_io_wt_actv_nz_0_14),
    .io_wt_actv_nz_0_15(u_active_io_wt_actv_nz_0_15),
    .io_wt_actv_nz_0_16(u_active_io_wt_actv_nz_0_16),
    .io_wt_actv_nz_0_17(u_active_io_wt_actv_nz_0_17),
    .io_wt_actv_nz_0_18(u_active_io_wt_actv_nz_0_18),
    .io_wt_actv_nz_0_19(u_active_io_wt_actv_nz_0_19),
    .io_wt_actv_nz_0_20(u_active_io_wt_actv_nz_0_20),
    .io_wt_actv_nz_0_21(u_active_io_wt_actv_nz_0_21),
    .io_wt_actv_nz_0_22(u_active_io_wt_actv_nz_0_22),
    .io_wt_actv_nz_0_23(u_active_io_wt_actv_nz_0_23),
    .io_wt_actv_nz_0_24(u_active_io_wt_actv_nz_0_24),
    .io_wt_actv_nz_0_25(u_active_io_wt_actv_nz_0_25),
    .io_wt_actv_nz_0_26(u_active_io_wt_actv_nz_0_26),
    .io_wt_actv_nz_0_27(u_active_io_wt_actv_nz_0_27),
    .io_wt_actv_nz_0_28(u_active_io_wt_actv_nz_0_28),
    .io_wt_actv_nz_0_29(u_active_io_wt_actv_nz_0_29),
    .io_wt_actv_nz_0_30(u_active_io_wt_actv_nz_0_30),
    .io_wt_actv_nz_0_31(u_active_io_wt_actv_nz_0_31),
    .io_wt_actv_nz_0_32(u_active_io_wt_actv_nz_0_32),
    .io_wt_actv_nz_0_33(u_active_io_wt_actv_nz_0_33),
    .io_wt_actv_nz_0_34(u_active_io_wt_actv_nz_0_34),
    .io_wt_actv_nz_0_35(u_active_io_wt_actv_nz_0_35),
    .io_wt_actv_nz_0_36(u_active_io_wt_actv_nz_0_36),
    .io_wt_actv_nz_0_37(u_active_io_wt_actv_nz_0_37),
    .io_wt_actv_nz_0_38(u_active_io_wt_actv_nz_0_38),
    .io_wt_actv_nz_0_39(u_active_io_wt_actv_nz_0_39),
    .io_wt_actv_nz_0_40(u_active_io_wt_actv_nz_0_40),
    .io_wt_actv_nz_0_41(u_active_io_wt_actv_nz_0_41),
    .io_wt_actv_nz_0_42(u_active_io_wt_actv_nz_0_42),
    .io_wt_actv_nz_0_43(u_active_io_wt_actv_nz_0_43),
    .io_wt_actv_nz_0_44(u_active_io_wt_actv_nz_0_44),
    .io_wt_actv_nz_0_45(u_active_io_wt_actv_nz_0_45),
    .io_wt_actv_nz_0_46(u_active_io_wt_actv_nz_0_46),
    .io_wt_actv_nz_0_47(u_active_io_wt_actv_nz_0_47),
    .io_wt_actv_nz_0_48(u_active_io_wt_actv_nz_0_48),
    .io_wt_actv_nz_0_49(u_active_io_wt_actv_nz_0_49),
    .io_wt_actv_nz_0_50(u_active_io_wt_actv_nz_0_50),
    .io_wt_actv_nz_0_51(u_active_io_wt_actv_nz_0_51),
    .io_wt_actv_nz_0_52(u_active_io_wt_actv_nz_0_52),
    .io_wt_actv_nz_0_53(u_active_io_wt_actv_nz_0_53),
    .io_wt_actv_nz_0_54(u_active_io_wt_actv_nz_0_54),
    .io_wt_actv_nz_0_55(u_active_io_wt_actv_nz_0_55),
    .io_wt_actv_nz_0_56(u_active_io_wt_actv_nz_0_56),
    .io_wt_actv_nz_0_57(u_active_io_wt_actv_nz_0_57),
    .io_wt_actv_nz_0_58(u_active_io_wt_actv_nz_0_58),
    .io_wt_actv_nz_0_59(u_active_io_wt_actv_nz_0_59),
    .io_wt_actv_nz_0_60(u_active_io_wt_actv_nz_0_60),
    .io_wt_actv_nz_0_61(u_active_io_wt_actv_nz_0_61),
    .io_wt_actv_nz_0_62(u_active_io_wt_actv_nz_0_62),
    .io_wt_actv_nz_0_63(u_active_io_wt_actv_nz_0_63),
    .io_wt_actv_nz_0_64(u_active_io_wt_actv_nz_0_64),
    .io_wt_actv_nz_0_65(u_active_io_wt_actv_nz_0_65),
    .io_wt_actv_nz_0_66(u_active_io_wt_actv_nz_0_66),
    .io_wt_actv_nz_0_67(u_active_io_wt_actv_nz_0_67),
    .io_wt_actv_nz_0_68(u_active_io_wt_actv_nz_0_68),
    .io_wt_actv_nz_0_69(u_active_io_wt_actv_nz_0_69),
    .io_wt_actv_nz_0_70(u_active_io_wt_actv_nz_0_70),
    .io_wt_actv_nz_0_71(u_active_io_wt_actv_nz_0_71),
    .io_wt_actv_nz_0_72(u_active_io_wt_actv_nz_0_72),
    .io_wt_actv_nz_0_73(u_active_io_wt_actv_nz_0_73),
    .io_wt_actv_nz_0_74(u_active_io_wt_actv_nz_0_74),
    .io_wt_actv_nz_0_75(u_active_io_wt_actv_nz_0_75),
    .io_wt_actv_nz_0_76(u_active_io_wt_actv_nz_0_76),
    .io_wt_actv_nz_0_77(u_active_io_wt_actv_nz_0_77),
    .io_wt_actv_nz_0_78(u_active_io_wt_actv_nz_0_78),
    .io_wt_actv_nz_0_79(u_active_io_wt_actv_nz_0_79),
    .io_wt_actv_nz_0_80(u_active_io_wt_actv_nz_0_80),
    .io_wt_actv_nz_0_81(u_active_io_wt_actv_nz_0_81),
    .io_wt_actv_nz_0_82(u_active_io_wt_actv_nz_0_82),
    .io_wt_actv_nz_0_83(u_active_io_wt_actv_nz_0_83),
    .io_wt_actv_nz_0_84(u_active_io_wt_actv_nz_0_84),
    .io_wt_actv_nz_0_85(u_active_io_wt_actv_nz_0_85),
    .io_wt_actv_nz_0_86(u_active_io_wt_actv_nz_0_86),
    .io_wt_actv_nz_0_87(u_active_io_wt_actv_nz_0_87),
    .io_wt_actv_nz_0_88(u_active_io_wt_actv_nz_0_88),
    .io_wt_actv_nz_0_89(u_active_io_wt_actv_nz_0_89),
    .io_wt_actv_nz_0_90(u_active_io_wt_actv_nz_0_90),
    .io_wt_actv_nz_0_91(u_active_io_wt_actv_nz_0_91),
    .io_wt_actv_nz_0_92(u_active_io_wt_actv_nz_0_92),
    .io_wt_actv_nz_0_93(u_active_io_wt_actv_nz_0_93),
    .io_wt_actv_nz_0_94(u_active_io_wt_actv_nz_0_94),
    .io_wt_actv_nz_0_95(u_active_io_wt_actv_nz_0_95),
    .io_wt_actv_nz_0_96(u_active_io_wt_actv_nz_0_96),
    .io_wt_actv_nz_0_97(u_active_io_wt_actv_nz_0_97),
    .io_wt_actv_nz_0_98(u_active_io_wt_actv_nz_0_98),
    .io_wt_actv_nz_0_99(u_active_io_wt_actv_nz_0_99),
    .io_wt_actv_nz_0_100(u_active_io_wt_actv_nz_0_100),
    .io_wt_actv_nz_0_101(u_active_io_wt_actv_nz_0_101),
    .io_wt_actv_nz_0_102(u_active_io_wt_actv_nz_0_102),
    .io_wt_actv_nz_0_103(u_active_io_wt_actv_nz_0_103),
    .io_wt_actv_nz_0_104(u_active_io_wt_actv_nz_0_104),
    .io_wt_actv_nz_0_105(u_active_io_wt_actv_nz_0_105),
    .io_wt_actv_nz_0_106(u_active_io_wt_actv_nz_0_106),
    .io_wt_actv_nz_0_107(u_active_io_wt_actv_nz_0_107),
    .io_wt_actv_nz_0_108(u_active_io_wt_actv_nz_0_108),
    .io_wt_actv_nz_0_109(u_active_io_wt_actv_nz_0_109),
    .io_wt_actv_nz_0_110(u_active_io_wt_actv_nz_0_110),
    .io_wt_actv_nz_0_111(u_active_io_wt_actv_nz_0_111),
    .io_wt_actv_nz_0_112(u_active_io_wt_actv_nz_0_112),
    .io_wt_actv_nz_0_113(u_active_io_wt_actv_nz_0_113),
    .io_wt_actv_nz_0_114(u_active_io_wt_actv_nz_0_114),
    .io_wt_actv_nz_0_115(u_active_io_wt_actv_nz_0_115),
    .io_wt_actv_nz_0_116(u_active_io_wt_actv_nz_0_116),
    .io_wt_actv_nz_0_117(u_active_io_wt_actv_nz_0_117),
    .io_wt_actv_nz_0_118(u_active_io_wt_actv_nz_0_118),
    .io_wt_actv_nz_0_119(u_active_io_wt_actv_nz_0_119),
    .io_wt_actv_nz_0_120(u_active_io_wt_actv_nz_0_120),
    .io_wt_actv_nz_0_121(u_active_io_wt_actv_nz_0_121),
    .io_wt_actv_nz_0_122(u_active_io_wt_actv_nz_0_122),
    .io_wt_actv_nz_0_123(u_active_io_wt_actv_nz_0_123),
    .io_wt_actv_nz_0_124(u_active_io_wt_actv_nz_0_124),
    .io_wt_actv_nz_0_125(u_active_io_wt_actv_nz_0_125),
    .io_wt_actv_nz_0_126(u_active_io_wt_actv_nz_0_126),
    .io_wt_actv_nz_0_127(u_active_io_wt_actv_nz_0_127),
    .io_wt_actv_pvld_0_0(u_active_io_wt_actv_pvld_0_0),
    .io_wt_actv_pvld_0_1(u_active_io_wt_actv_pvld_0_1),
    .io_wt_actv_pvld_0_2(u_active_io_wt_actv_pvld_0_2),
    .io_wt_actv_pvld_0_3(u_active_io_wt_actv_pvld_0_3),
    .io_wt_actv_pvld_0_4(u_active_io_wt_actv_pvld_0_4),
    .io_wt_actv_pvld_0_5(u_active_io_wt_actv_pvld_0_5),
    .io_wt_actv_pvld_0_6(u_active_io_wt_actv_pvld_0_6),
    .io_wt_actv_pvld_0_7(u_active_io_wt_actv_pvld_0_7),
    .io_wt_actv_pvld_0_8(u_active_io_wt_actv_pvld_0_8),
    .io_wt_actv_pvld_0_9(u_active_io_wt_actv_pvld_0_9),
    .io_wt_actv_pvld_0_10(u_active_io_wt_actv_pvld_0_10),
    .io_wt_actv_pvld_0_11(u_active_io_wt_actv_pvld_0_11),
    .io_wt_actv_pvld_0_12(u_active_io_wt_actv_pvld_0_12),
    .io_wt_actv_pvld_0_13(u_active_io_wt_actv_pvld_0_13),
    .io_wt_actv_pvld_0_14(u_active_io_wt_actv_pvld_0_14),
    .io_wt_actv_pvld_0_15(u_active_io_wt_actv_pvld_0_15),
    .io_wt_actv_pvld_0_16(u_active_io_wt_actv_pvld_0_16),
    .io_wt_actv_pvld_0_17(u_active_io_wt_actv_pvld_0_17),
    .io_wt_actv_pvld_0_18(u_active_io_wt_actv_pvld_0_18),
    .io_wt_actv_pvld_0_19(u_active_io_wt_actv_pvld_0_19),
    .io_wt_actv_pvld_0_20(u_active_io_wt_actv_pvld_0_20),
    .io_wt_actv_pvld_0_21(u_active_io_wt_actv_pvld_0_21),
    .io_wt_actv_pvld_0_22(u_active_io_wt_actv_pvld_0_22),
    .io_wt_actv_pvld_0_23(u_active_io_wt_actv_pvld_0_23),
    .io_wt_actv_pvld_0_24(u_active_io_wt_actv_pvld_0_24),
    .io_wt_actv_pvld_0_25(u_active_io_wt_actv_pvld_0_25),
    .io_wt_actv_pvld_0_26(u_active_io_wt_actv_pvld_0_26),
    .io_wt_actv_pvld_0_27(u_active_io_wt_actv_pvld_0_27),
    .io_wt_actv_pvld_0_28(u_active_io_wt_actv_pvld_0_28),
    .io_wt_actv_pvld_0_29(u_active_io_wt_actv_pvld_0_29),
    .io_wt_actv_pvld_0_30(u_active_io_wt_actv_pvld_0_30),
    .io_wt_actv_pvld_0_31(u_active_io_wt_actv_pvld_0_31),
    .io_wt_actv_pvld_0_32(u_active_io_wt_actv_pvld_0_32),
    .io_wt_actv_pvld_0_33(u_active_io_wt_actv_pvld_0_33),
    .io_wt_actv_pvld_0_34(u_active_io_wt_actv_pvld_0_34),
    .io_wt_actv_pvld_0_35(u_active_io_wt_actv_pvld_0_35),
    .io_wt_actv_pvld_0_36(u_active_io_wt_actv_pvld_0_36),
    .io_wt_actv_pvld_0_37(u_active_io_wt_actv_pvld_0_37),
    .io_wt_actv_pvld_0_38(u_active_io_wt_actv_pvld_0_38),
    .io_wt_actv_pvld_0_39(u_active_io_wt_actv_pvld_0_39),
    .io_wt_actv_pvld_0_40(u_active_io_wt_actv_pvld_0_40),
    .io_wt_actv_pvld_0_41(u_active_io_wt_actv_pvld_0_41),
    .io_wt_actv_pvld_0_42(u_active_io_wt_actv_pvld_0_42),
    .io_wt_actv_pvld_0_43(u_active_io_wt_actv_pvld_0_43),
    .io_wt_actv_pvld_0_44(u_active_io_wt_actv_pvld_0_44),
    .io_wt_actv_pvld_0_45(u_active_io_wt_actv_pvld_0_45),
    .io_wt_actv_pvld_0_46(u_active_io_wt_actv_pvld_0_46),
    .io_wt_actv_pvld_0_47(u_active_io_wt_actv_pvld_0_47),
    .io_wt_actv_pvld_0_48(u_active_io_wt_actv_pvld_0_48),
    .io_wt_actv_pvld_0_49(u_active_io_wt_actv_pvld_0_49),
    .io_wt_actv_pvld_0_50(u_active_io_wt_actv_pvld_0_50),
    .io_wt_actv_pvld_0_51(u_active_io_wt_actv_pvld_0_51),
    .io_wt_actv_pvld_0_52(u_active_io_wt_actv_pvld_0_52),
    .io_wt_actv_pvld_0_53(u_active_io_wt_actv_pvld_0_53),
    .io_wt_actv_pvld_0_54(u_active_io_wt_actv_pvld_0_54),
    .io_wt_actv_pvld_0_55(u_active_io_wt_actv_pvld_0_55),
    .io_wt_actv_pvld_0_56(u_active_io_wt_actv_pvld_0_56),
    .io_wt_actv_pvld_0_57(u_active_io_wt_actv_pvld_0_57),
    .io_wt_actv_pvld_0_58(u_active_io_wt_actv_pvld_0_58),
    .io_wt_actv_pvld_0_59(u_active_io_wt_actv_pvld_0_59),
    .io_wt_actv_pvld_0_60(u_active_io_wt_actv_pvld_0_60),
    .io_wt_actv_pvld_0_61(u_active_io_wt_actv_pvld_0_61),
    .io_wt_actv_pvld_0_62(u_active_io_wt_actv_pvld_0_62),
    .io_wt_actv_pvld_0_63(u_active_io_wt_actv_pvld_0_63),
    .io_wt_actv_pvld_0_64(u_active_io_wt_actv_pvld_0_64),
    .io_wt_actv_pvld_0_65(u_active_io_wt_actv_pvld_0_65),
    .io_wt_actv_pvld_0_66(u_active_io_wt_actv_pvld_0_66),
    .io_wt_actv_pvld_0_67(u_active_io_wt_actv_pvld_0_67),
    .io_wt_actv_pvld_0_68(u_active_io_wt_actv_pvld_0_68),
    .io_wt_actv_pvld_0_69(u_active_io_wt_actv_pvld_0_69),
    .io_wt_actv_pvld_0_70(u_active_io_wt_actv_pvld_0_70),
    .io_wt_actv_pvld_0_71(u_active_io_wt_actv_pvld_0_71),
    .io_wt_actv_pvld_0_72(u_active_io_wt_actv_pvld_0_72),
    .io_wt_actv_pvld_0_73(u_active_io_wt_actv_pvld_0_73),
    .io_wt_actv_pvld_0_74(u_active_io_wt_actv_pvld_0_74),
    .io_wt_actv_pvld_0_75(u_active_io_wt_actv_pvld_0_75),
    .io_wt_actv_pvld_0_76(u_active_io_wt_actv_pvld_0_76),
    .io_wt_actv_pvld_0_77(u_active_io_wt_actv_pvld_0_77),
    .io_wt_actv_pvld_0_78(u_active_io_wt_actv_pvld_0_78),
    .io_wt_actv_pvld_0_79(u_active_io_wt_actv_pvld_0_79),
    .io_wt_actv_pvld_0_80(u_active_io_wt_actv_pvld_0_80),
    .io_wt_actv_pvld_0_81(u_active_io_wt_actv_pvld_0_81),
    .io_wt_actv_pvld_0_82(u_active_io_wt_actv_pvld_0_82),
    .io_wt_actv_pvld_0_83(u_active_io_wt_actv_pvld_0_83),
    .io_wt_actv_pvld_0_84(u_active_io_wt_actv_pvld_0_84),
    .io_wt_actv_pvld_0_85(u_active_io_wt_actv_pvld_0_85),
    .io_wt_actv_pvld_0_86(u_active_io_wt_actv_pvld_0_86),
    .io_wt_actv_pvld_0_87(u_active_io_wt_actv_pvld_0_87),
    .io_wt_actv_pvld_0_88(u_active_io_wt_actv_pvld_0_88),
    .io_wt_actv_pvld_0_89(u_active_io_wt_actv_pvld_0_89),
    .io_wt_actv_pvld_0_90(u_active_io_wt_actv_pvld_0_90),
    .io_wt_actv_pvld_0_91(u_active_io_wt_actv_pvld_0_91),
    .io_wt_actv_pvld_0_92(u_active_io_wt_actv_pvld_0_92),
    .io_wt_actv_pvld_0_93(u_active_io_wt_actv_pvld_0_93),
    .io_wt_actv_pvld_0_94(u_active_io_wt_actv_pvld_0_94),
    .io_wt_actv_pvld_0_95(u_active_io_wt_actv_pvld_0_95),
    .io_wt_actv_pvld_0_96(u_active_io_wt_actv_pvld_0_96),
    .io_wt_actv_pvld_0_97(u_active_io_wt_actv_pvld_0_97),
    .io_wt_actv_pvld_0_98(u_active_io_wt_actv_pvld_0_98),
    .io_wt_actv_pvld_0_99(u_active_io_wt_actv_pvld_0_99),
    .io_wt_actv_pvld_0_100(u_active_io_wt_actv_pvld_0_100),
    .io_wt_actv_pvld_0_101(u_active_io_wt_actv_pvld_0_101),
    .io_wt_actv_pvld_0_102(u_active_io_wt_actv_pvld_0_102),
    .io_wt_actv_pvld_0_103(u_active_io_wt_actv_pvld_0_103),
    .io_wt_actv_pvld_0_104(u_active_io_wt_actv_pvld_0_104),
    .io_wt_actv_pvld_0_105(u_active_io_wt_actv_pvld_0_105),
    .io_wt_actv_pvld_0_106(u_active_io_wt_actv_pvld_0_106),
    .io_wt_actv_pvld_0_107(u_active_io_wt_actv_pvld_0_107),
    .io_wt_actv_pvld_0_108(u_active_io_wt_actv_pvld_0_108),
    .io_wt_actv_pvld_0_109(u_active_io_wt_actv_pvld_0_109),
    .io_wt_actv_pvld_0_110(u_active_io_wt_actv_pvld_0_110),
    .io_wt_actv_pvld_0_111(u_active_io_wt_actv_pvld_0_111),
    .io_wt_actv_pvld_0_112(u_active_io_wt_actv_pvld_0_112),
    .io_wt_actv_pvld_0_113(u_active_io_wt_actv_pvld_0_113),
    .io_wt_actv_pvld_0_114(u_active_io_wt_actv_pvld_0_114),
    .io_wt_actv_pvld_0_115(u_active_io_wt_actv_pvld_0_115),
    .io_wt_actv_pvld_0_116(u_active_io_wt_actv_pvld_0_116),
    .io_wt_actv_pvld_0_117(u_active_io_wt_actv_pvld_0_117),
    .io_wt_actv_pvld_0_118(u_active_io_wt_actv_pvld_0_118),
    .io_wt_actv_pvld_0_119(u_active_io_wt_actv_pvld_0_119),
    .io_wt_actv_pvld_0_120(u_active_io_wt_actv_pvld_0_120),
    .io_wt_actv_pvld_0_121(u_active_io_wt_actv_pvld_0_121),
    .io_wt_actv_pvld_0_122(u_active_io_wt_actv_pvld_0_122),
    .io_wt_actv_pvld_0_123(u_active_io_wt_actv_pvld_0_123),
    .io_wt_actv_pvld_0_124(u_active_io_wt_actv_pvld_0_124),
    .io_wt_actv_pvld_0_125(u_active_io_wt_actv_pvld_0_125),
    .io_wt_actv_pvld_0_126(u_active_io_wt_actv_pvld_0_126),
    .io_wt_actv_pvld_0_127(u_active_io_wt_actv_pvld_0_127)
  );
  NV_NVDLA_CMAC_CORE_mac NV_NVDLA_CMAC_CORE_mac ( // @[NV_NVDLA_CMAC_core.scala 108:56]
    .clock(NV_NVDLA_CMAC_CORE_mac_clock),
    .io_dat_actv_data_0(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_0),
    .io_dat_actv_data_1(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_1),
    .io_dat_actv_data_2(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_2),
    .io_dat_actv_data_3(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_3),
    .io_dat_actv_data_4(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_4),
    .io_dat_actv_data_5(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_5),
    .io_dat_actv_data_6(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_6),
    .io_dat_actv_data_7(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_7),
    .io_dat_actv_data_8(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_8),
    .io_dat_actv_data_9(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_9),
    .io_dat_actv_data_10(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_10),
    .io_dat_actv_data_11(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_11),
    .io_dat_actv_data_12(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_12),
    .io_dat_actv_data_13(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_13),
    .io_dat_actv_data_14(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_14),
    .io_dat_actv_data_15(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_15),
    .io_dat_actv_data_16(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_16),
    .io_dat_actv_data_17(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_17),
    .io_dat_actv_data_18(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_18),
    .io_dat_actv_data_19(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_19),
    .io_dat_actv_data_20(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_20),
    .io_dat_actv_data_21(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_21),
    .io_dat_actv_data_22(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_22),
    .io_dat_actv_data_23(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_23),
    .io_dat_actv_data_24(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_24),
    .io_dat_actv_data_25(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_25),
    .io_dat_actv_data_26(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_26),
    .io_dat_actv_data_27(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_27),
    .io_dat_actv_data_28(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_28),
    .io_dat_actv_data_29(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_29),
    .io_dat_actv_data_30(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_30),
    .io_dat_actv_data_31(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_31),
    .io_dat_actv_data_32(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_32),
    .io_dat_actv_data_33(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_33),
    .io_dat_actv_data_34(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_34),
    .io_dat_actv_data_35(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_35),
    .io_dat_actv_data_36(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_36),
    .io_dat_actv_data_37(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_37),
    .io_dat_actv_data_38(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_38),
    .io_dat_actv_data_39(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_39),
    .io_dat_actv_data_40(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_40),
    .io_dat_actv_data_41(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_41),
    .io_dat_actv_data_42(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_42),
    .io_dat_actv_data_43(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_43),
    .io_dat_actv_data_44(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_44),
    .io_dat_actv_data_45(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_45),
    .io_dat_actv_data_46(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_46),
    .io_dat_actv_data_47(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_47),
    .io_dat_actv_data_48(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_48),
    .io_dat_actv_data_49(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_49),
    .io_dat_actv_data_50(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_50),
    .io_dat_actv_data_51(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_51),
    .io_dat_actv_data_52(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_52),
    .io_dat_actv_data_53(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_53),
    .io_dat_actv_data_54(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_54),
    .io_dat_actv_data_55(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_55),
    .io_dat_actv_data_56(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_56),
    .io_dat_actv_data_57(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_57),
    .io_dat_actv_data_58(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_58),
    .io_dat_actv_data_59(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_59),
    .io_dat_actv_data_60(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_60),
    .io_dat_actv_data_61(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_61),
    .io_dat_actv_data_62(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_62),
    .io_dat_actv_data_63(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_63),
    .io_dat_actv_data_64(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_64),
    .io_dat_actv_data_65(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_65),
    .io_dat_actv_data_66(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_66),
    .io_dat_actv_data_67(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_67),
    .io_dat_actv_data_68(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_68),
    .io_dat_actv_data_69(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_69),
    .io_dat_actv_data_70(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_70),
    .io_dat_actv_data_71(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_71),
    .io_dat_actv_data_72(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_72),
    .io_dat_actv_data_73(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_73),
    .io_dat_actv_data_74(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_74),
    .io_dat_actv_data_75(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_75),
    .io_dat_actv_data_76(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_76),
    .io_dat_actv_data_77(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_77),
    .io_dat_actv_data_78(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_78),
    .io_dat_actv_data_79(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_79),
    .io_dat_actv_data_80(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_80),
    .io_dat_actv_data_81(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_81),
    .io_dat_actv_data_82(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_82),
    .io_dat_actv_data_83(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_83),
    .io_dat_actv_data_84(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_84),
    .io_dat_actv_data_85(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_85),
    .io_dat_actv_data_86(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_86),
    .io_dat_actv_data_87(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_87),
    .io_dat_actv_data_88(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_88),
    .io_dat_actv_data_89(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_89),
    .io_dat_actv_data_90(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_90),
    .io_dat_actv_data_91(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_91),
    .io_dat_actv_data_92(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_92),
    .io_dat_actv_data_93(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_93),
    .io_dat_actv_data_94(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_94),
    .io_dat_actv_data_95(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_95),
    .io_dat_actv_data_96(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_96),
    .io_dat_actv_data_97(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_97),
    .io_dat_actv_data_98(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_98),
    .io_dat_actv_data_99(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_99),
    .io_dat_actv_data_100(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_100),
    .io_dat_actv_data_101(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_101),
    .io_dat_actv_data_102(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_102),
    .io_dat_actv_data_103(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_103),
    .io_dat_actv_data_104(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_104),
    .io_dat_actv_data_105(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_105),
    .io_dat_actv_data_106(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_106),
    .io_dat_actv_data_107(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_107),
    .io_dat_actv_data_108(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_108),
    .io_dat_actv_data_109(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_109),
    .io_dat_actv_data_110(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_110),
    .io_dat_actv_data_111(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_111),
    .io_dat_actv_data_112(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_112),
    .io_dat_actv_data_113(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_113),
    .io_dat_actv_data_114(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_114),
    .io_dat_actv_data_115(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_115),
    .io_dat_actv_data_116(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_116),
    .io_dat_actv_data_117(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_117),
    .io_dat_actv_data_118(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_118),
    .io_dat_actv_data_119(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_119),
    .io_dat_actv_data_120(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_120),
    .io_dat_actv_data_121(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_121),
    .io_dat_actv_data_122(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_122),
    .io_dat_actv_data_123(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_123),
    .io_dat_actv_data_124(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_124),
    .io_dat_actv_data_125(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_125),
    .io_dat_actv_data_126(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_126),
    .io_dat_actv_data_127(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_127),
    .io_dat_actv_nz_0(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_0),
    .io_dat_actv_nz_1(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_1),
    .io_dat_actv_nz_2(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_2),
    .io_dat_actv_nz_3(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_3),
    .io_dat_actv_nz_4(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_4),
    .io_dat_actv_nz_5(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_5),
    .io_dat_actv_nz_6(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_6),
    .io_dat_actv_nz_7(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_7),
    .io_dat_actv_nz_8(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_8),
    .io_dat_actv_nz_9(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_9),
    .io_dat_actv_nz_10(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_10),
    .io_dat_actv_nz_11(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_11),
    .io_dat_actv_nz_12(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_12),
    .io_dat_actv_nz_13(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_13),
    .io_dat_actv_nz_14(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_14),
    .io_dat_actv_nz_15(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_15),
    .io_dat_actv_nz_16(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_16),
    .io_dat_actv_nz_17(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_17),
    .io_dat_actv_nz_18(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_18),
    .io_dat_actv_nz_19(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_19),
    .io_dat_actv_nz_20(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_20),
    .io_dat_actv_nz_21(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_21),
    .io_dat_actv_nz_22(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_22),
    .io_dat_actv_nz_23(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_23),
    .io_dat_actv_nz_24(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_24),
    .io_dat_actv_nz_25(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_25),
    .io_dat_actv_nz_26(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_26),
    .io_dat_actv_nz_27(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_27),
    .io_dat_actv_nz_28(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_28),
    .io_dat_actv_nz_29(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_29),
    .io_dat_actv_nz_30(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_30),
    .io_dat_actv_nz_31(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_31),
    .io_dat_actv_nz_32(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_32),
    .io_dat_actv_nz_33(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_33),
    .io_dat_actv_nz_34(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_34),
    .io_dat_actv_nz_35(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_35),
    .io_dat_actv_nz_36(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_36),
    .io_dat_actv_nz_37(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_37),
    .io_dat_actv_nz_38(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_38),
    .io_dat_actv_nz_39(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_39),
    .io_dat_actv_nz_40(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_40),
    .io_dat_actv_nz_41(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_41),
    .io_dat_actv_nz_42(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_42),
    .io_dat_actv_nz_43(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_43),
    .io_dat_actv_nz_44(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_44),
    .io_dat_actv_nz_45(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_45),
    .io_dat_actv_nz_46(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_46),
    .io_dat_actv_nz_47(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_47),
    .io_dat_actv_nz_48(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_48),
    .io_dat_actv_nz_49(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_49),
    .io_dat_actv_nz_50(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_50),
    .io_dat_actv_nz_51(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_51),
    .io_dat_actv_nz_52(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_52),
    .io_dat_actv_nz_53(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_53),
    .io_dat_actv_nz_54(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_54),
    .io_dat_actv_nz_55(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_55),
    .io_dat_actv_nz_56(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_56),
    .io_dat_actv_nz_57(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_57),
    .io_dat_actv_nz_58(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_58),
    .io_dat_actv_nz_59(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_59),
    .io_dat_actv_nz_60(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_60),
    .io_dat_actv_nz_61(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_61),
    .io_dat_actv_nz_62(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_62),
    .io_dat_actv_nz_63(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_63),
    .io_dat_actv_nz_64(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_64),
    .io_dat_actv_nz_65(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_65),
    .io_dat_actv_nz_66(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_66),
    .io_dat_actv_nz_67(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_67),
    .io_dat_actv_nz_68(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_68),
    .io_dat_actv_nz_69(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_69),
    .io_dat_actv_nz_70(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_70),
    .io_dat_actv_nz_71(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_71),
    .io_dat_actv_nz_72(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_72),
    .io_dat_actv_nz_73(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_73),
    .io_dat_actv_nz_74(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_74),
    .io_dat_actv_nz_75(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_75),
    .io_dat_actv_nz_76(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_76),
    .io_dat_actv_nz_77(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_77),
    .io_dat_actv_nz_78(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_78),
    .io_dat_actv_nz_79(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_79),
    .io_dat_actv_nz_80(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_80),
    .io_dat_actv_nz_81(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_81),
    .io_dat_actv_nz_82(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_82),
    .io_dat_actv_nz_83(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_83),
    .io_dat_actv_nz_84(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_84),
    .io_dat_actv_nz_85(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_85),
    .io_dat_actv_nz_86(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_86),
    .io_dat_actv_nz_87(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_87),
    .io_dat_actv_nz_88(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_88),
    .io_dat_actv_nz_89(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_89),
    .io_dat_actv_nz_90(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_90),
    .io_dat_actv_nz_91(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_91),
    .io_dat_actv_nz_92(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_92),
    .io_dat_actv_nz_93(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_93),
    .io_dat_actv_nz_94(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_94),
    .io_dat_actv_nz_95(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_95),
    .io_dat_actv_nz_96(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_96),
    .io_dat_actv_nz_97(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_97),
    .io_dat_actv_nz_98(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_98),
    .io_dat_actv_nz_99(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_99),
    .io_dat_actv_nz_100(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_100),
    .io_dat_actv_nz_101(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_101),
    .io_dat_actv_nz_102(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_102),
    .io_dat_actv_nz_103(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_103),
    .io_dat_actv_nz_104(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_104),
    .io_dat_actv_nz_105(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_105),
    .io_dat_actv_nz_106(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_106),
    .io_dat_actv_nz_107(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_107),
    .io_dat_actv_nz_108(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_108),
    .io_dat_actv_nz_109(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_109),
    .io_dat_actv_nz_110(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_110),
    .io_dat_actv_nz_111(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_111),
    .io_dat_actv_nz_112(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_112),
    .io_dat_actv_nz_113(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_113),
    .io_dat_actv_nz_114(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_114),
    .io_dat_actv_nz_115(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_115),
    .io_dat_actv_nz_116(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_116),
    .io_dat_actv_nz_117(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_117),
    .io_dat_actv_nz_118(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_118),
    .io_dat_actv_nz_119(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_119),
    .io_dat_actv_nz_120(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_120),
    .io_dat_actv_nz_121(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_121),
    .io_dat_actv_nz_122(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_122),
    .io_dat_actv_nz_123(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_123),
    .io_dat_actv_nz_124(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_124),
    .io_dat_actv_nz_125(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_125),
    .io_dat_actv_nz_126(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_126),
    .io_dat_actv_nz_127(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_127),
    .io_dat_actv_pvld_0(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_0),
    .io_dat_actv_pvld_1(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_1),
    .io_dat_actv_pvld_2(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_2),
    .io_dat_actv_pvld_3(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_3),
    .io_dat_actv_pvld_4(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_4),
    .io_dat_actv_pvld_5(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_5),
    .io_dat_actv_pvld_6(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_6),
    .io_dat_actv_pvld_7(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_7),
    .io_dat_actv_pvld_8(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_8),
    .io_dat_actv_pvld_9(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_9),
    .io_dat_actv_pvld_10(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_10),
    .io_dat_actv_pvld_11(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_11),
    .io_dat_actv_pvld_12(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_12),
    .io_dat_actv_pvld_13(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_13),
    .io_dat_actv_pvld_14(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_14),
    .io_dat_actv_pvld_15(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_15),
    .io_dat_actv_pvld_16(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_16),
    .io_dat_actv_pvld_17(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_17),
    .io_dat_actv_pvld_18(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_18),
    .io_dat_actv_pvld_19(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_19),
    .io_dat_actv_pvld_20(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_20),
    .io_dat_actv_pvld_21(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_21),
    .io_dat_actv_pvld_22(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_22),
    .io_dat_actv_pvld_23(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_23),
    .io_dat_actv_pvld_24(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_24),
    .io_dat_actv_pvld_25(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_25),
    .io_dat_actv_pvld_26(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_26),
    .io_dat_actv_pvld_27(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_27),
    .io_dat_actv_pvld_28(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_28),
    .io_dat_actv_pvld_29(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_29),
    .io_dat_actv_pvld_30(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_30),
    .io_dat_actv_pvld_31(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_31),
    .io_dat_actv_pvld_32(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_32),
    .io_dat_actv_pvld_33(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_33),
    .io_dat_actv_pvld_34(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_34),
    .io_dat_actv_pvld_35(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_35),
    .io_dat_actv_pvld_36(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_36),
    .io_dat_actv_pvld_37(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_37),
    .io_dat_actv_pvld_38(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_38),
    .io_dat_actv_pvld_39(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_39),
    .io_dat_actv_pvld_40(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_40),
    .io_dat_actv_pvld_41(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_41),
    .io_dat_actv_pvld_42(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_42),
    .io_dat_actv_pvld_43(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_43),
    .io_dat_actv_pvld_44(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_44),
    .io_dat_actv_pvld_45(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_45),
    .io_dat_actv_pvld_46(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_46),
    .io_dat_actv_pvld_47(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_47),
    .io_dat_actv_pvld_48(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_48),
    .io_dat_actv_pvld_49(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_49),
    .io_dat_actv_pvld_50(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_50),
    .io_dat_actv_pvld_51(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_51),
    .io_dat_actv_pvld_52(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_52),
    .io_dat_actv_pvld_53(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_53),
    .io_dat_actv_pvld_54(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_54),
    .io_dat_actv_pvld_55(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_55),
    .io_dat_actv_pvld_56(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_56),
    .io_dat_actv_pvld_57(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_57),
    .io_dat_actv_pvld_58(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_58),
    .io_dat_actv_pvld_59(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_59),
    .io_dat_actv_pvld_60(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_60),
    .io_dat_actv_pvld_61(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_61),
    .io_dat_actv_pvld_62(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_62),
    .io_dat_actv_pvld_63(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_63),
    .io_dat_actv_pvld_64(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_64),
    .io_dat_actv_pvld_65(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_65),
    .io_dat_actv_pvld_66(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_66),
    .io_dat_actv_pvld_67(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_67),
    .io_dat_actv_pvld_68(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_68),
    .io_dat_actv_pvld_69(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_69),
    .io_dat_actv_pvld_70(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_70),
    .io_dat_actv_pvld_71(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_71),
    .io_dat_actv_pvld_72(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_72),
    .io_dat_actv_pvld_73(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_73),
    .io_dat_actv_pvld_74(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_74),
    .io_dat_actv_pvld_75(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_75),
    .io_dat_actv_pvld_76(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_76),
    .io_dat_actv_pvld_77(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_77),
    .io_dat_actv_pvld_78(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_78),
    .io_dat_actv_pvld_79(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_79),
    .io_dat_actv_pvld_80(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_80),
    .io_dat_actv_pvld_81(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_81),
    .io_dat_actv_pvld_82(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_82),
    .io_dat_actv_pvld_83(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_83),
    .io_dat_actv_pvld_84(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_84),
    .io_dat_actv_pvld_85(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_85),
    .io_dat_actv_pvld_86(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_86),
    .io_dat_actv_pvld_87(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_87),
    .io_dat_actv_pvld_88(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_88),
    .io_dat_actv_pvld_89(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_89),
    .io_dat_actv_pvld_90(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_90),
    .io_dat_actv_pvld_91(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_91),
    .io_dat_actv_pvld_92(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_92),
    .io_dat_actv_pvld_93(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_93),
    .io_dat_actv_pvld_94(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_94),
    .io_dat_actv_pvld_95(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_95),
    .io_dat_actv_pvld_96(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_96),
    .io_dat_actv_pvld_97(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_97),
    .io_dat_actv_pvld_98(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_98),
    .io_dat_actv_pvld_99(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_99),
    .io_dat_actv_pvld_100(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_100),
    .io_dat_actv_pvld_101(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_101),
    .io_dat_actv_pvld_102(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_102),
    .io_dat_actv_pvld_103(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_103),
    .io_dat_actv_pvld_104(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_104),
    .io_dat_actv_pvld_105(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_105),
    .io_dat_actv_pvld_106(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_106),
    .io_dat_actv_pvld_107(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_107),
    .io_dat_actv_pvld_108(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_108),
    .io_dat_actv_pvld_109(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_109),
    .io_dat_actv_pvld_110(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_110),
    .io_dat_actv_pvld_111(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_111),
    .io_dat_actv_pvld_112(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_112),
    .io_dat_actv_pvld_113(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_113),
    .io_dat_actv_pvld_114(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_114),
    .io_dat_actv_pvld_115(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_115),
    .io_dat_actv_pvld_116(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_116),
    .io_dat_actv_pvld_117(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_117),
    .io_dat_actv_pvld_118(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_118),
    .io_dat_actv_pvld_119(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_119),
    .io_dat_actv_pvld_120(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_120),
    .io_dat_actv_pvld_121(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_121),
    .io_dat_actv_pvld_122(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_122),
    .io_dat_actv_pvld_123(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_123),
    .io_dat_actv_pvld_124(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_124),
    .io_dat_actv_pvld_125(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_125),
    .io_dat_actv_pvld_126(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_126),
    .io_dat_actv_pvld_127(NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_127),
    .io_wt_actv_data_0(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_0),
    .io_wt_actv_data_1(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_1),
    .io_wt_actv_data_2(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_2),
    .io_wt_actv_data_3(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_3),
    .io_wt_actv_data_4(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_4),
    .io_wt_actv_data_5(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_5),
    .io_wt_actv_data_6(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_6),
    .io_wt_actv_data_7(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_7),
    .io_wt_actv_data_8(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_8),
    .io_wt_actv_data_9(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_9),
    .io_wt_actv_data_10(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_10),
    .io_wt_actv_data_11(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_11),
    .io_wt_actv_data_12(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_12),
    .io_wt_actv_data_13(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_13),
    .io_wt_actv_data_14(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_14),
    .io_wt_actv_data_15(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_15),
    .io_wt_actv_data_16(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_16),
    .io_wt_actv_data_17(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_17),
    .io_wt_actv_data_18(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_18),
    .io_wt_actv_data_19(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_19),
    .io_wt_actv_data_20(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_20),
    .io_wt_actv_data_21(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_21),
    .io_wt_actv_data_22(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_22),
    .io_wt_actv_data_23(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_23),
    .io_wt_actv_data_24(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_24),
    .io_wt_actv_data_25(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_25),
    .io_wt_actv_data_26(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_26),
    .io_wt_actv_data_27(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_27),
    .io_wt_actv_data_28(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_28),
    .io_wt_actv_data_29(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_29),
    .io_wt_actv_data_30(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_30),
    .io_wt_actv_data_31(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_31),
    .io_wt_actv_data_32(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_32),
    .io_wt_actv_data_33(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_33),
    .io_wt_actv_data_34(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_34),
    .io_wt_actv_data_35(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_35),
    .io_wt_actv_data_36(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_36),
    .io_wt_actv_data_37(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_37),
    .io_wt_actv_data_38(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_38),
    .io_wt_actv_data_39(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_39),
    .io_wt_actv_data_40(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_40),
    .io_wt_actv_data_41(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_41),
    .io_wt_actv_data_42(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_42),
    .io_wt_actv_data_43(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_43),
    .io_wt_actv_data_44(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_44),
    .io_wt_actv_data_45(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_45),
    .io_wt_actv_data_46(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_46),
    .io_wt_actv_data_47(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_47),
    .io_wt_actv_data_48(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_48),
    .io_wt_actv_data_49(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_49),
    .io_wt_actv_data_50(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_50),
    .io_wt_actv_data_51(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_51),
    .io_wt_actv_data_52(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_52),
    .io_wt_actv_data_53(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_53),
    .io_wt_actv_data_54(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_54),
    .io_wt_actv_data_55(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_55),
    .io_wt_actv_data_56(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_56),
    .io_wt_actv_data_57(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_57),
    .io_wt_actv_data_58(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_58),
    .io_wt_actv_data_59(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_59),
    .io_wt_actv_data_60(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_60),
    .io_wt_actv_data_61(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_61),
    .io_wt_actv_data_62(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_62),
    .io_wt_actv_data_63(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_63),
    .io_wt_actv_data_64(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_64),
    .io_wt_actv_data_65(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_65),
    .io_wt_actv_data_66(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_66),
    .io_wt_actv_data_67(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_67),
    .io_wt_actv_data_68(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_68),
    .io_wt_actv_data_69(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_69),
    .io_wt_actv_data_70(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_70),
    .io_wt_actv_data_71(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_71),
    .io_wt_actv_data_72(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_72),
    .io_wt_actv_data_73(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_73),
    .io_wt_actv_data_74(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_74),
    .io_wt_actv_data_75(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_75),
    .io_wt_actv_data_76(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_76),
    .io_wt_actv_data_77(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_77),
    .io_wt_actv_data_78(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_78),
    .io_wt_actv_data_79(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_79),
    .io_wt_actv_data_80(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_80),
    .io_wt_actv_data_81(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_81),
    .io_wt_actv_data_82(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_82),
    .io_wt_actv_data_83(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_83),
    .io_wt_actv_data_84(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_84),
    .io_wt_actv_data_85(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_85),
    .io_wt_actv_data_86(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_86),
    .io_wt_actv_data_87(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_87),
    .io_wt_actv_data_88(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_88),
    .io_wt_actv_data_89(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_89),
    .io_wt_actv_data_90(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_90),
    .io_wt_actv_data_91(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_91),
    .io_wt_actv_data_92(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_92),
    .io_wt_actv_data_93(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_93),
    .io_wt_actv_data_94(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_94),
    .io_wt_actv_data_95(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_95),
    .io_wt_actv_data_96(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_96),
    .io_wt_actv_data_97(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_97),
    .io_wt_actv_data_98(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_98),
    .io_wt_actv_data_99(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_99),
    .io_wt_actv_data_100(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_100),
    .io_wt_actv_data_101(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_101),
    .io_wt_actv_data_102(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_102),
    .io_wt_actv_data_103(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_103),
    .io_wt_actv_data_104(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_104),
    .io_wt_actv_data_105(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_105),
    .io_wt_actv_data_106(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_106),
    .io_wt_actv_data_107(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_107),
    .io_wt_actv_data_108(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_108),
    .io_wt_actv_data_109(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_109),
    .io_wt_actv_data_110(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_110),
    .io_wt_actv_data_111(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_111),
    .io_wt_actv_data_112(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_112),
    .io_wt_actv_data_113(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_113),
    .io_wt_actv_data_114(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_114),
    .io_wt_actv_data_115(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_115),
    .io_wt_actv_data_116(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_116),
    .io_wt_actv_data_117(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_117),
    .io_wt_actv_data_118(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_118),
    .io_wt_actv_data_119(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_119),
    .io_wt_actv_data_120(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_120),
    .io_wt_actv_data_121(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_121),
    .io_wt_actv_data_122(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_122),
    .io_wt_actv_data_123(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_123),
    .io_wt_actv_data_124(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_124),
    .io_wt_actv_data_125(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_125),
    .io_wt_actv_data_126(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_126),
    .io_wt_actv_data_127(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_127),
    .io_wt_actv_nz_0(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_0),
    .io_wt_actv_nz_1(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_1),
    .io_wt_actv_nz_2(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_2),
    .io_wt_actv_nz_3(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_3),
    .io_wt_actv_nz_4(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_4),
    .io_wt_actv_nz_5(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_5),
    .io_wt_actv_nz_6(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_6),
    .io_wt_actv_nz_7(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_7),
    .io_wt_actv_nz_8(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_8),
    .io_wt_actv_nz_9(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_9),
    .io_wt_actv_nz_10(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_10),
    .io_wt_actv_nz_11(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_11),
    .io_wt_actv_nz_12(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_12),
    .io_wt_actv_nz_13(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_13),
    .io_wt_actv_nz_14(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_14),
    .io_wt_actv_nz_15(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_15),
    .io_wt_actv_nz_16(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_16),
    .io_wt_actv_nz_17(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_17),
    .io_wt_actv_nz_18(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_18),
    .io_wt_actv_nz_19(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_19),
    .io_wt_actv_nz_20(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_20),
    .io_wt_actv_nz_21(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_21),
    .io_wt_actv_nz_22(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_22),
    .io_wt_actv_nz_23(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_23),
    .io_wt_actv_nz_24(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_24),
    .io_wt_actv_nz_25(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_25),
    .io_wt_actv_nz_26(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_26),
    .io_wt_actv_nz_27(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_27),
    .io_wt_actv_nz_28(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_28),
    .io_wt_actv_nz_29(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_29),
    .io_wt_actv_nz_30(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_30),
    .io_wt_actv_nz_31(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_31),
    .io_wt_actv_nz_32(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_32),
    .io_wt_actv_nz_33(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_33),
    .io_wt_actv_nz_34(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_34),
    .io_wt_actv_nz_35(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_35),
    .io_wt_actv_nz_36(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_36),
    .io_wt_actv_nz_37(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_37),
    .io_wt_actv_nz_38(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_38),
    .io_wt_actv_nz_39(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_39),
    .io_wt_actv_nz_40(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_40),
    .io_wt_actv_nz_41(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_41),
    .io_wt_actv_nz_42(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_42),
    .io_wt_actv_nz_43(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_43),
    .io_wt_actv_nz_44(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_44),
    .io_wt_actv_nz_45(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_45),
    .io_wt_actv_nz_46(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_46),
    .io_wt_actv_nz_47(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_47),
    .io_wt_actv_nz_48(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_48),
    .io_wt_actv_nz_49(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_49),
    .io_wt_actv_nz_50(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_50),
    .io_wt_actv_nz_51(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_51),
    .io_wt_actv_nz_52(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_52),
    .io_wt_actv_nz_53(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_53),
    .io_wt_actv_nz_54(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_54),
    .io_wt_actv_nz_55(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_55),
    .io_wt_actv_nz_56(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_56),
    .io_wt_actv_nz_57(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_57),
    .io_wt_actv_nz_58(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_58),
    .io_wt_actv_nz_59(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_59),
    .io_wt_actv_nz_60(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_60),
    .io_wt_actv_nz_61(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_61),
    .io_wt_actv_nz_62(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_62),
    .io_wt_actv_nz_63(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_63),
    .io_wt_actv_nz_64(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_64),
    .io_wt_actv_nz_65(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_65),
    .io_wt_actv_nz_66(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_66),
    .io_wt_actv_nz_67(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_67),
    .io_wt_actv_nz_68(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_68),
    .io_wt_actv_nz_69(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_69),
    .io_wt_actv_nz_70(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_70),
    .io_wt_actv_nz_71(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_71),
    .io_wt_actv_nz_72(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_72),
    .io_wt_actv_nz_73(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_73),
    .io_wt_actv_nz_74(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_74),
    .io_wt_actv_nz_75(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_75),
    .io_wt_actv_nz_76(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_76),
    .io_wt_actv_nz_77(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_77),
    .io_wt_actv_nz_78(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_78),
    .io_wt_actv_nz_79(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_79),
    .io_wt_actv_nz_80(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_80),
    .io_wt_actv_nz_81(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_81),
    .io_wt_actv_nz_82(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_82),
    .io_wt_actv_nz_83(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_83),
    .io_wt_actv_nz_84(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_84),
    .io_wt_actv_nz_85(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_85),
    .io_wt_actv_nz_86(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_86),
    .io_wt_actv_nz_87(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_87),
    .io_wt_actv_nz_88(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_88),
    .io_wt_actv_nz_89(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_89),
    .io_wt_actv_nz_90(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_90),
    .io_wt_actv_nz_91(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_91),
    .io_wt_actv_nz_92(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_92),
    .io_wt_actv_nz_93(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_93),
    .io_wt_actv_nz_94(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_94),
    .io_wt_actv_nz_95(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_95),
    .io_wt_actv_nz_96(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_96),
    .io_wt_actv_nz_97(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_97),
    .io_wt_actv_nz_98(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_98),
    .io_wt_actv_nz_99(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_99),
    .io_wt_actv_nz_100(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_100),
    .io_wt_actv_nz_101(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_101),
    .io_wt_actv_nz_102(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_102),
    .io_wt_actv_nz_103(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_103),
    .io_wt_actv_nz_104(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_104),
    .io_wt_actv_nz_105(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_105),
    .io_wt_actv_nz_106(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_106),
    .io_wt_actv_nz_107(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_107),
    .io_wt_actv_nz_108(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_108),
    .io_wt_actv_nz_109(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_109),
    .io_wt_actv_nz_110(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_110),
    .io_wt_actv_nz_111(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_111),
    .io_wt_actv_nz_112(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_112),
    .io_wt_actv_nz_113(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_113),
    .io_wt_actv_nz_114(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_114),
    .io_wt_actv_nz_115(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_115),
    .io_wt_actv_nz_116(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_116),
    .io_wt_actv_nz_117(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_117),
    .io_wt_actv_nz_118(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_118),
    .io_wt_actv_nz_119(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_119),
    .io_wt_actv_nz_120(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_120),
    .io_wt_actv_nz_121(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_121),
    .io_wt_actv_nz_122(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_122),
    .io_wt_actv_nz_123(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_123),
    .io_wt_actv_nz_124(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_124),
    .io_wt_actv_nz_125(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_125),
    .io_wt_actv_nz_126(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_126),
    .io_wt_actv_nz_127(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_127),
    .io_wt_actv_pvld_0(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_0),
    .io_wt_actv_pvld_1(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_1),
    .io_wt_actv_pvld_2(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_2),
    .io_wt_actv_pvld_3(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_3),
    .io_wt_actv_pvld_4(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_4),
    .io_wt_actv_pvld_5(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_5),
    .io_wt_actv_pvld_6(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_6),
    .io_wt_actv_pvld_7(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_7),
    .io_wt_actv_pvld_8(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_8),
    .io_wt_actv_pvld_9(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_9),
    .io_wt_actv_pvld_10(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_10),
    .io_wt_actv_pvld_11(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_11),
    .io_wt_actv_pvld_12(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_12),
    .io_wt_actv_pvld_13(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_13),
    .io_wt_actv_pvld_14(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_14),
    .io_wt_actv_pvld_15(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_15),
    .io_wt_actv_pvld_16(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_16),
    .io_wt_actv_pvld_17(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_17),
    .io_wt_actv_pvld_18(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_18),
    .io_wt_actv_pvld_19(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_19),
    .io_wt_actv_pvld_20(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_20),
    .io_wt_actv_pvld_21(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_21),
    .io_wt_actv_pvld_22(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_22),
    .io_wt_actv_pvld_23(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_23),
    .io_wt_actv_pvld_24(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_24),
    .io_wt_actv_pvld_25(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_25),
    .io_wt_actv_pvld_26(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_26),
    .io_wt_actv_pvld_27(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_27),
    .io_wt_actv_pvld_28(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_28),
    .io_wt_actv_pvld_29(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_29),
    .io_wt_actv_pvld_30(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_30),
    .io_wt_actv_pvld_31(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_31),
    .io_wt_actv_pvld_32(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_32),
    .io_wt_actv_pvld_33(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_33),
    .io_wt_actv_pvld_34(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_34),
    .io_wt_actv_pvld_35(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_35),
    .io_wt_actv_pvld_36(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_36),
    .io_wt_actv_pvld_37(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_37),
    .io_wt_actv_pvld_38(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_38),
    .io_wt_actv_pvld_39(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_39),
    .io_wt_actv_pvld_40(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_40),
    .io_wt_actv_pvld_41(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_41),
    .io_wt_actv_pvld_42(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_42),
    .io_wt_actv_pvld_43(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_43),
    .io_wt_actv_pvld_44(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_44),
    .io_wt_actv_pvld_45(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_45),
    .io_wt_actv_pvld_46(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_46),
    .io_wt_actv_pvld_47(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_47),
    .io_wt_actv_pvld_48(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_48),
    .io_wt_actv_pvld_49(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_49),
    .io_wt_actv_pvld_50(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_50),
    .io_wt_actv_pvld_51(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_51),
    .io_wt_actv_pvld_52(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_52),
    .io_wt_actv_pvld_53(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_53),
    .io_wt_actv_pvld_54(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_54),
    .io_wt_actv_pvld_55(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_55),
    .io_wt_actv_pvld_56(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_56),
    .io_wt_actv_pvld_57(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_57),
    .io_wt_actv_pvld_58(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_58),
    .io_wt_actv_pvld_59(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_59),
    .io_wt_actv_pvld_60(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_60),
    .io_wt_actv_pvld_61(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_61),
    .io_wt_actv_pvld_62(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_62),
    .io_wt_actv_pvld_63(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_63),
    .io_wt_actv_pvld_64(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_64),
    .io_wt_actv_pvld_65(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_65),
    .io_wt_actv_pvld_66(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_66),
    .io_wt_actv_pvld_67(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_67),
    .io_wt_actv_pvld_68(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_68),
    .io_wt_actv_pvld_69(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_69),
    .io_wt_actv_pvld_70(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_70),
    .io_wt_actv_pvld_71(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_71),
    .io_wt_actv_pvld_72(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_72),
    .io_wt_actv_pvld_73(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_73),
    .io_wt_actv_pvld_74(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_74),
    .io_wt_actv_pvld_75(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_75),
    .io_wt_actv_pvld_76(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_76),
    .io_wt_actv_pvld_77(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_77),
    .io_wt_actv_pvld_78(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_78),
    .io_wt_actv_pvld_79(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_79),
    .io_wt_actv_pvld_80(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_80),
    .io_wt_actv_pvld_81(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_81),
    .io_wt_actv_pvld_82(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_82),
    .io_wt_actv_pvld_83(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_83),
    .io_wt_actv_pvld_84(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_84),
    .io_wt_actv_pvld_85(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_85),
    .io_wt_actv_pvld_86(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_86),
    .io_wt_actv_pvld_87(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_87),
    .io_wt_actv_pvld_88(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_88),
    .io_wt_actv_pvld_89(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_89),
    .io_wt_actv_pvld_90(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_90),
    .io_wt_actv_pvld_91(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_91),
    .io_wt_actv_pvld_92(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_92),
    .io_wt_actv_pvld_93(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_93),
    .io_wt_actv_pvld_94(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_94),
    .io_wt_actv_pvld_95(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_95),
    .io_wt_actv_pvld_96(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_96),
    .io_wt_actv_pvld_97(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_97),
    .io_wt_actv_pvld_98(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_98),
    .io_wt_actv_pvld_99(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_99),
    .io_wt_actv_pvld_100(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_100),
    .io_wt_actv_pvld_101(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_101),
    .io_wt_actv_pvld_102(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_102),
    .io_wt_actv_pvld_103(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_103),
    .io_wt_actv_pvld_104(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_104),
    .io_wt_actv_pvld_105(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_105),
    .io_wt_actv_pvld_106(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_106),
    .io_wt_actv_pvld_107(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_107),
    .io_wt_actv_pvld_108(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_108),
    .io_wt_actv_pvld_109(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_109),
    .io_wt_actv_pvld_110(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_110),
    .io_wt_actv_pvld_111(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_111),
    .io_wt_actv_pvld_112(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_112),
    .io_wt_actv_pvld_113(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_113),
    .io_wt_actv_pvld_114(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_114),
    .io_wt_actv_pvld_115(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_115),
    .io_wt_actv_pvld_116(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_116),
    .io_wt_actv_pvld_117(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_117),
    .io_wt_actv_pvld_118(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_118),
    .io_wt_actv_pvld_119(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_119),
    .io_wt_actv_pvld_120(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_120),
    .io_wt_actv_pvld_121(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_121),
    .io_wt_actv_pvld_122(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_122),
    .io_wt_actv_pvld_123(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_123),
    .io_wt_actv_pvld_124(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_124),
    .io_wt_actv_pvld_125(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_125),
    .io_wt_actv_pvld_126(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_126),
    .io_wt_actv_pvld_127(NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_127),
    .io_mac_out_data(NV_NVDLA_CMAC_CORE_mac_io_mac_out_data),
    .io_mac_out_pvld(NV_NVDLA_CMAC_CORE_mac_io_mac_out_pvld)
  );
  NV_NVDLA_CMAC_CORE_rt_out u_rt_out ( // @[NV_NVDLA_CMAC_core.scala 129:26]
    .clock(u_rt_out_clock),
    .reset(u_rt_out_reset),
    .io_out_data_0(u_rt_out_io_out_data_0),
    .io_out_mask_0(u_rt_out_io_out_mask_0),
    .io_out_pd(u_rt_out_io_out_pd),
    .io_out_pvld(u_rt_out_io_out_pvld),
    .io_mac2accu_data_0(u_rt_out_io_mac2accu_data_0),
    .io_mac2accu_mask_0(u_rt_out_io_mac2accu_mask_0),
    .io_mac2accu_pd(u_rt_out_io_mac2accu_pd),
    .io_mac2accu_pvld(u_rt_out_io_mac2accu_pvld),
    .io_dp2reg_done(u_rt_out_io_dp2reg_done)
  );
  assign io_mac2accu_pvld = u_rt_out_io_mac2accu_pvld; // @[NV_NVDLA_CMAC_core.scala 140:22]
  assign io_mac2accu_mask_0 = u_rt_out_io_mac2accu_mask_0; // @[NV_NVDLA_CMAC_core.scala 138:22]
  assign io_mac2accu_data_0 = u_rt_out_io_mac2accu_data_0; // @[NV_NVDLA_CMAC_core.scala 137:22]
  assign io_mac2accu_pd = u_rt_out_io_mac2accu_pd; // @[NV_NVDLA_CMAC_core.scala 139:20]
  assign io_dp2reg_done = u_rt_out_io_dp2reg_done; // @[NV_NVDLA_CMAC_core.scala 136:20]
  assign u_rt_in_clock = clock;
  assign u_rt_in_reset = reset;
  assign u_rt_in_io_sc2mac_dat_data_0 = io_sc2mac_dat_data_0; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_1 = io_sc2mac_dat_data_1; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_2 = io_sc2mac_dat_data_2; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_3 = io_sc2mac_dat_data_3; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_4 = io_sc2mac_dat_data_4; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_5 = io_sc2mac_dat_data_5; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_6 = io_sc2mac_dat_data_6; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_7 = io_sc2mac_dat_data_7; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_8 = io_sc2mac_dat_data_8; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_9 = io_sc2mac_dat_data_9; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_10 = io_sc2mac_dat_data_10; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_11 = io_sc2mac_dat_data_11; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_12 = io_sc2mac_dat_data_12; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_13 = io_sc2mac_dat_data_13; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_14 = io_sc2mac_dat_data_14; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_15 = io_sc2mac_dat_data_15; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_16 = io_sc2mac_dat_data_16; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_17 = io_sc2mac_dat_data_17; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_18 = io_sc2mac_dat_data_18; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_19 = io_sc2mac_dat_data_19; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_20 = io_sc2mac_dat_data_20; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_21 = io_sc2mac_dat_data_21; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_22 = io_sc2mac_dat_data_22; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_23 = io_sc2mac_dat_data_23; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_24 = io_sc2mac_dat_data_24; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_25 = io_sc2mac_dat_data_25; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_26 = io_sc2mac_dat_data_26; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_27 = io_sc2mac_dat_data_27; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_28 = io_sc2mac_dat_data_28; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_29 = io_sc2mac_dat_data_29; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_30 = io_sc2mac_dat_data_30; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_31 = io_sc2mac_dat_data_31; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_32 = io_sc2mac_dat_data_32; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_33 = io_sc2mac_dat_data_33; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_34 = io_sc2mac_dat_data_34; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_35 = io_sc2mac_dat_data_35; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_36 = io_sc2mac_dat_data_36; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_37 = io_sc2mac_dat_data_37; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_38 = io_sc2mac_dat_data_38; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_39 = io_sc2mac_dat_data_39; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_40 = io_sc2mac_dat_data_40; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_41 = io_sc2mac_dat_data_41; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_42 = io_sc2mac_dat_data_42; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_43 = io_sc2mac_dat_data_43; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_44 = io_sc2mac_dat_data_44; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_45 = io_sc2mac_dat_data_45; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_46 = io_sc2mac_dat_data_46; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_47 = io_sc2mac_dat_data_47; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_48 = io_sc2mac_dat_data_48; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_49 = io_sc2mac_dat_data_49; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_50 = io_sc2mac_dat_data_50; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_51 = io_sc2mac_dat_data_51; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_52 = io_sc2mac_dat_data_52; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_53 = io_sc2mac_dat_data_53; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_54 = io_sc2mac_dat_data_54; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_55 = io_sc2mac_dat_data_55; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_56 = io_sc2mac_dat_data_56; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_57 = io_sc2mac_dat_data_57; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_58 = io_sc2mac_dat_data_58; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_59 = io_sc2mac_dat_data_59; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_60 = io_sc2mac_dat_data_60; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_61 = io_sc2mac_dat_data_61; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_62 = io_sc2mac_dat_data_62; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_63 = io_sc2mac_dat_data_63; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_64 = io_sc2mac_dat_data_64; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_65 = io_sc2mac_dat_data_65; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_66 = io_sc2mac_dat_data_66; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_67 = io_sc2mac_dat_data_67; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_68 = io_sc2mac_dat_data_68; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_69 = io_sc2mac_dat_data_69; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_70 = io_sc2mac_dat_data_70; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_71 = io_sc2mac_dat_data_71; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_72 = io_sc2mac_dat_data_72; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_73 = io_sc2mac_dat_data_73; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_74 = io_sc2mac_dat_data_74; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_75 = io_sc2mac_dat_data_75; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_76 = io_sc2mac_dat_data_76; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_77 = io_sc2mac_dat_data_77; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_78 = io_sc2mac_dat_data_78; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_79 = io_sc2mac_dat_data_79; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_80 = io_sc2mac_dat_data_80; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_81 = io_sc2mac_dat_data_81; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_82 = io_sc2mac_dat_data_82; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_83 = io_sc2mac_dat_data_83; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_84 = io_sc2mac_dat_data_84; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_85 = io_sc2mac_dat_data_85; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_86 = io_sc2mac_dat_data_86; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_87 = io_sc2mac_dat_data_87; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_88 = io_sc2mac_dat_data_88; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_89 = io_sc2mac_dat_data_89; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_90 = io_sc2mac_dat_data_90; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_91 = io_sc2mac_dat_data_91; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_92 = io_sc2mac_dat_data_92; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_93 = io_sc2mac_dat_data_93; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_94 = io_sc2mac_dat_data_94; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_95 = io_sc2mac_dat_data_95; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_96 = io_sc2mac_dat_data_96; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_97 = io_sc2mac_dat_data_97; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_98 = io_sc2mac_dat_data_98; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_99 = io_sc2mac_dat_data_99; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_100 = io_sc2mac_dat_data_100; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_101 = io_sc2mac_dat_data_101; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_102 = io_sc2mac_dat_data_102; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_103 = io_sc2mac_dat_data_103; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_104 = io_sc2mac_dat_data_104; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_105 = io_sc2mac_dat_data_105; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_106 = io_sc2mac_dat_data_106; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_107 = io_sc2mac_dat_data_107; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_108 = io_sc2mac_dat_data_108; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_109 = io_sc2mac_dat_data_109; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_110 = io_sc2mac_dat_data_110; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_111 = io_sc2mac_dat_data_111; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_112 = io_sc2mac_dat_data_112; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_113 = io_sc2mac_dat_data_113; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_114 = io_sc2mac_dat_data_114; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_115 = io_sc2mac_dat_data_115; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_116 = io_sc2mac_dat_data_116; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_117 = io_sc2mac_dat_data_117; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_118 = io_sc2mac_dat_data_118; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_119 = io_sc2mac_dat_data_119; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_120 = io_sc2mac_dat_data_120; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_121 = io_sc2mac_dat_data_121; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_122 = io_sc2mac_dat_data_122; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_123 = io_sc2mac_dat_data_123; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_124 = io_sc2mac_dat_data_124; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_125 = io_sc2mac_dat_data_125; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_126 = io_sc2mac_dat_data_126; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_data_127 = io_sc2mac_dat_data_127; // @[NV_NVDLA_CMAC_core.scala 56:32]
  assign u_rt_in_io_sc2mac_dat_mask_0 = io_sc2mac_dat_mask_0; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_1 = io_sc2mac_dat_mask_1; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_2 = io_sc2mac_dat_mask_2; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_3 = io_sc2mac_dat_mask_3; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_4 = io_sc2mac_dat_mask_4; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_5 = io_sc2mac_dat_mask_5; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_6 = io_sc2mac_dat_mask_6; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_7 = io_sc2mac_dat_mask_7; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_8 = io_sc2mac_dat_mask_8; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_9 = io_sc2mac_dat_mask_9; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_10 = io_sc2mac_dat_mask_10; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_11 = io_sc2mac_dat_mask_11; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_12 = io_sc2mac_dat_mask_12; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_13 = io_sc2mac_dat_mask_13; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_14 = io_sc2mac_dat_mask_14; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_15 = io_sc2mac_dat_mask_15; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_16 = io_sc2mac_dat_mask_16; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_17 = io_sc2mac_dat_mask_17; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_18 = io_sc2mac_dat_mask_18; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_19 = io_sc2mac_dat_mask_19; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_20 = io_sc2mac_dat_mask_20; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_21 = io_sc2mac_dat_mask_21; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_22 = io_sc2mac_dat_mask_22; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_23 = io_sc2mac_dat_mask_23; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_24 = io_sc2mac_dat_mask_24; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_25 = io_sc2mac_dat_mask_25; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_26 = io_sc2mac_dat_mask_26; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_27 = io_sc2mac_dat_mask_27; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_28 = io_sc2mac_dat_mask_28; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_29 = io_sc2mac_dat_mask_29; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_30 = io_sc2mac_dat_mask_30; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_31 = io_sc2mac_dat_mask_31; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_32 = io_sc2mac_dat_mask_32; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_33 = io_sc2mac_dat_mask_33; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_34 = io_sc2mac_dat_mask_34; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_35 = io_sc2mac_dat_mask_35; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_36 = io_sc2mac_dat_mask_36; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_37 = io_sc2mac_dat_mask_37; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_38 = io_sc2mac_dat_mask_38; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_39 = io_sc2mac_dat_mask_39; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_40 = io_sc2mac_dat_mask_40; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_41 = io_sc2mac_dat_mask_41; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_42 = io_sc2mac_dat_mask_42; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_43 = io_sc2mac_dat_mask_43; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_44 = io_sc2mac_dat_mask_44; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_45 = io_sc2mac_dat_mask_45; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_46 = io_sc2mac_dat_mask_46; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_47 = io_sc2mac_dat_mask_47; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_48 = io_sc2mac_dat_mask_48; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_49 = io_sc2mac_dat_mask_49; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_50 = io_sc2mac_dat_mask_50; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_51 = io_sc2mac_dat_mask_51; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_52 = io_sc2mac_dat_mask_52; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_53 = io_sc2mac_dat_mask_53; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_54 = io_sc2mac_dat_mask_54; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_55 = io_sc2mac_dat_mask_55; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_56 = io_sc2mac_dat_mask_56; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_57 = io_sc2mac_dat_mask_57; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_58 = io_sc2mac_dat_mask_58; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_59 = io_sc2mac_dat_mask_59; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_60 = io_sc2mac_dat_mask_60; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_61 = io_sc2mac_dat_mask_61; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_62 = io_sc2mac_dat_mask_62; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_63 = io_sc2mac_dat_mask_63; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_64 = io_sc2mac_dat_mask_64; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_65 = io_sc2mac_dat_mask_65; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_66 = io_sc2mac_dat_mask_66; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_67 = io_sc2mac_dat_mask_67; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_68 = io_sc2mac_dat_mask_68; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_69 = io_sc2mac_dat_mask_69; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_70 = io_sc2mac_dat_mask_70; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_71 = io_sc2mac_dat_mask_71; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_72 = io_sc2mac_dat_mask_72; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_73 = io_sc2mac_dat_mask_73; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_74 = io_sc2mac_dat_mask_74; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_75 = io_sc2mac_dat_mask_75; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_76 = io_sc2mac_dat_mask_76; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_77 = io_sc2mac_dat_mask_77; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_78 = io_sc2mac_dat_mask_78; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_79 = io_sc2mac_dat_mask_79; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_80 = io_sc2mac_dat_mask_80; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_81 = io_sc2mac_dat_mask_81; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_82 = io_sc2mac_dat_mask_82; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_83 = io_sc2mac_dat_mask_83; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_84 = io_sc2mac_dat_mask_84; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_85 = io_sc2mac_dat_mask_85; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_86 = io_sc2mac_dat_mask_86; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_87 = io_sc2mac_dat_mask_87; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_88 = io_sc2mac_dat_mask_88; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_89 = io_sc2mac_dat_mask_89; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_90 = io_sc2mac_dat_mask_90; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_91 = io_sc2mac_dat_mask_91; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_92 = io_sc2mac_dat_mask_92; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_93 = io_sc2mac_dat_mask_93; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_94 = io_sc2mac_dat_mask_94; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_95 = io_sc2mac_dat_mask_95; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_96 = io_sc2mac_dat_mask_96; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_97 = io_sc2mac_dat_mask_97; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_98 = io_sc2mac_dat_mask_98; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_99 = io_sc2mac_dat_mask_99; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_100 = io_sc2mac_dat_mask_100; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_101 = io_sc2mac_dat_mask_101; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_102 = io_sc2mac_dat_mask_102; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_103 = io_sc2mac_dat_mask_103; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_104 = io_sc2mac_dat_mask_104; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_105 = io_sc2mac_dat_mask_105; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_106 = io_sc2mac_dat_mask_106; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_107 = io_sc2mac_dat_mask_107; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_108 = io_sc2mac_dat_mask_108; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_109 = io_sc2mac_dat_mask_109; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_110 = io_sc2mac_dat_mask_110; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_111 = io_sc2mac_dat_mask_111; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_112 = io_sc2mac_dat_mask_112; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_113 = io_sc2mac_dat_mask_113; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_114 = io_sc2mac_dat_mask_114; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_115 = io_sc2mac_dat_mask_115; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_116 = io_sc2mac_dat_mask_116; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_117 = io_sc2mac_dat_mask_117; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_118 = io_sc2mac_dat_mask_118; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_119 = io_sc2mac_dat_mask_119; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_120 = io_sc2mac_dat_mask_120; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_121 = io_sc2mac_dat_mask_121; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_122 = io_sc2mac_dat_mask_122; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_123 = io_sc2mac_dat_mask_123; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_124 = io_sc2mac_dat_mask_124; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_125 = io_sc2mac_dat_mask_125; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_126 = io_sc2mac_dat_mask_126; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_mask_127 = io_sc2mac_dat_mask_127; // @[NV_NVDLA_CMAC_core.scala 55:32]
  assign u_rt_in_io_sc2mac_dat_pd = io_sc2mac_dat_pd; // @[NV_NVDLA_CMAC_core.scala 57:30]
  assign u_rt_in_io_sc2mac_dat_pvld = io_sc2mac_dat_pvld; // @[NV_NVDLA_CMAC_core.scala 54:32]
  assign u_rt_in_io_sc2mac_wt_data_0 = io_sc2mac_wt_data_0; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_1 = io_sc2mac_wt_data_1; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_2 = io_sc2mac_wt_data_2; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_3 = io_sc2mac_wt_data_3; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_4 = io_sc2mac_wt_data_4; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_5 = io_sc2mac_wt_data_5; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_6 = io_sc2mac_wt_data_6; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_7 = io_sc2mac_wt_data_7; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_8 = io_sc2mac_wt_data_8; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_9 = io_sc2mac_wt_data_9; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_10 = io_sc2mac_wt_data_10; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_11 = io_sc2mac_wt_data_11; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_12 = io_sc2mac_wt_data_12; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_13 = io_sc2mac_wt_data_13; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_14 = io_sc2mac_wt_data_14; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_15 = io_sc2mac_wt_data_15; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_16 = io_sc2mac_wt_data_16; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_17 = io_sc2mac_wt_data_17; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_18 = io_sc2mac_wt_data_18; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_19 = io_sc2mac_wt_data_19; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_20 = io_sc2mac_wt_data_20; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_21 = io_sc2mac_wt_data_21; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_22 = io_sc2mac_wt_data_22; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_23 = io_sc2mac_wt_data_23; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_24 = io_sc2mac_wt_data_24; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_25 = io_sc2mac_wt_data_25; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_26 = io_sc2mac_wt_data_26; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_27 = io_sc2mac_wt_data_27; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_28 = io_sc2mac_wt_data_28; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_29 = io_sc2mac_wt_data_29; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_30 = io_sc2mac_wt_data_30; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_31 = io_sc2mac_wt_data_31; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_32 = io_sc2mac_wt_data_32; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_33 = io_sc2mac_wt_data_33; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_34 = io_sc2mac_wt_data_34; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_35 = io_sc2mac_wt_data_35; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_36 = io_sc2mac_wt_data_36; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_37 = io_sc2mac_wt_data_37; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_38 = io_sc2mac_wt_data_38; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_39 = io_sc2mac_wt_data_39; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_40 = io_sc2mac_wt_data_40; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_41 = io_sc2mac_wt_data_41; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_42 = io_sc2mac_wt_data_42; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_43 = io_sc2mac_wt_data_43; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_44 = io_sc2mac_wt_data_44; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_45 = io_sc2mac_wt_data_45; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_46 = io_sc2mac_wt_data_46; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_47 = io_sc2mac_wt_data_47; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_48 = io_sc2mac_wt_data_48; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_49 = io_sc2mac_wt_data_49; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_50 = io_sc2mac_wt_data_50; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_51 = io_sc2mac_wt_data_51; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_52 = io_sc2mac_wt_data_52; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_53 = io_sc2mac_wt_data_53; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_54 = io_sc2mac_wt_data_54; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_55 = io_sc2mac_wt_data_55; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_56 = io_sc2mac_wt_data_56; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_57 = io_sc2mac_wt_data_57; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_58 = io_sc2mac_wt_data_58; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_59 = io_sc2mac_wt_data_59; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_60 = io_sc2mac_wt_data_60; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_61 = io_sc2mac_wt_data_61; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_62 = io_sc2mac_wt_data_62; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_63 = io_sc2mac_wt_data_63; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_64 = io_sc2mac_wt_data_64; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_65 = io_sc2mac_wt_data_65; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_66 = io_sc2mac_wt_data_66; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_67 = io_sc2mac_wt_data_67; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_68 = io_sc2mac_wt_data_68; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_69 = io_sc2mac_wt_data_69; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_70 = io_sc2mac_wt_data_70; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_71 = io_sc2mac_wt_data_71; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_72 = io_sc2mac_wt_data_72; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_73 = io_sc2mac_wt_data_73; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_74 = io_sc2mac_wt_data_74; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_75 = io_sc2mac_wt_data_75; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_76 = io_sc2mac_wt_data_76; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_77 = io_sc2mac_wt_data_77; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_78 = io_sc2mac_wt_data_78; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_79 = io_sc2mac_wt_data_79; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_80 = io_sc2mac_wt_data_80; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_81 = io_sc2mac_wt_data_81; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_82 = io_sc2mac_wt_data_82; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_83 = io_sc2mac_wt_data_83; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_84 = io_sc2mac_wt_data_84; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_85 = io_sc2mac_wt_data_85; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_86 = io_sc2mac_wt_data_86; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_87 = io_sc2mac_wt_data_87; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_88 = io_sc2mac_wt_data_88; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_89 = io_sc2mac_wt_data_89; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_90 = io_sc2mac_wt_data_90; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_91 = io_sc2mac_wt_data_91; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_92 = io_sc2mac_wt_data_92; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_93 = io_sc2mac_wt_data_93; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_94 = io_sc2mac_wt_data_94; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_95 = io_sc2mac_wt_data_95; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_96 = io_sc2mac_wt_data_96; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_97 = io_sc2mac_wt_data_97; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_98 = io_sc2mac_wt_data_98; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_99 = io_sc2mac_wt_data_99; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_100 = io_sc2mac_wt_data_100; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_101 = io_sc2mac_wt_data_101; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_102 = io_sc2mac_wt_data_102; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_103 = io_sc2mac_wt_data_103; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_104 = io_sc2mac_wt_data_104; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_105 = io_sc2mac_wt_data_105; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_106 = io_sc2mac_wt_data_106; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_107 = io_sc2mac_wt_data_107; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_108 = io_sc2mac_wt_data_108; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_109 = io_sc2mac_wt_data_109; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_110 = io_sc2mac_wt_data_110; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_111 = io_sc2mac_wt_data_111; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_112 = io_sc2mac_wt_data_112; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_113 = io_sc2mac_wt_data_113; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_114 = io_sc2mac_wt_data_114; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_115 = io_sc2mac_wt_data_115; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_116 = io_sc2mac_wt_data_116; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_117 = io_sc2mac_wt_data_117; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_118 = io_sc2mac_wt_data_118; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_119 = io_sc2mac_wt_data_119; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_120 = io_sc2mac_wt_data_120; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_121 = io_sc2mac_wt_data_121; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_122 = io_sc2mac_wt_data_122; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_123 = io_sc2mac_wt_data_123; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_124 = io_sc2mac_wt_data_124; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_125 = io_sc2mac_wt_data_125; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_126 = io_sc2mac_wt_data_126; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_data_127 = io_sc2mac_wt_data_127; // @[NV_NVDLA_CMAC_core.scala 61:31]
  assign u_rt_in_io_sc2mac_wt_mask_0 = io_sc2mac_wt_mask_0; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_1 = io_sc2mac_wt_mask_1; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_2 = io_sc2mac_wt_mask_2; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_3 = io_sc2mac_wt_mask_3; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_4 = io_sc2mac_wt_mask_4; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_5 = io_sc2mac_wt_mask_5; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_6 = io_sc2mac_wt_mask_6; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_7 = io_sc2mac_wt_mask_7; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_8 = io_sc2mac_wt_mask_8; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_9 = io_sc2mac_wt_mask_9; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_10 = io_sc2mac_wt_mask_10; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_11 = io_sc2mac_wt_mask_11; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_12 = io_sc2mac_wt_mask_12; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_13 = io_sc2mac_wt_mask_13; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_14 = io_sc2mac_wt_mask_14; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_15 = io_sc2mac_wt_mask_15; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_16 = io_sc2mac_wt_mask_16; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_17 = io_sc2mac_wt_mask_17; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_18 = io_sc2mac_wt_mask_18; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_19 = io_sc2mac_wt_mask_19; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_20 = io_sc2mac_wt_mask_20; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_21 = io_sc2mac_wt_mask_21; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_22 = io_sc2mac_wt_mask_22; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_23 = io_sc2mac_wt_mask_23; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_24 = io_sc2mac_wt_mask_24; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_25 = io_sc2mac_wt_mask_25; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_26 = io_sc2mac_wt_mask_26; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_27 = io_sc2mac_wt_mask_27; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_28 = io_sc2mac_wt_mask_28; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_29 = io_sc2mac_wt_mask_29; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_30 = io_sc2mac_wt_mask_30; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_31 = io_sc2mac_wt_mask_31; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_32 = io_sc2mac_wt_mask_32; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_33 = io_sc2mac_wt_mask_33; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_34 = io_sc2mac_wt_mask_34; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_35 = io_sc2mac_wt_mask_35; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_36 = io_sc2mac_wt_mask_36; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_37 = io_sc2mac_wt_mask_37; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_38 = io_sc2mac_wt_mask_38; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_39 = io_sc2mac_wt_mask_39; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_40 = io_sc2mac_wt_mask_40; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_41 = io_sc2mac_wt_mask_41; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_42 = io_sc2mac_wt_mask_42; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_43 = io_sc2mac_wt_mask_43; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_44 = io_sc2mac_wt_mask_44; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_45 = io_sc2mac_wt_mask_45; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_46 = io_sc2mac_wt_mask_46; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_47 = io_sc2mac_wt_mask_47; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_48 = io_sc2mac_wt_mask_48; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_49 = io_sc2mac_wt_mask_49; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_50 = io_sc2mac_wt_mask_50; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_51 = io_sc2mac_wt_mask_51; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_52 = io_sc2mac_wt_mask_52; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_53 = io_sc2mac_wt_mask_53; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_54 = io_sc2mac_wt_mask_54; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_55 = io_sc2mac_wt_mask_55; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_56 = io_sc2mac_wt_mask_56; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_57 = io_sc2mac_wt_mask_57; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_58 = io_sc2mac_wt_mask_58; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_59 = io_sc2mac_wt_mask_59; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_60 = io_sc2mac_wt_mask_60; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_61 = io_sc2mac_wt_mask_61; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_62 = io_sc2mac_wt_mask_62; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_63 = io_sc2mac_wt_mask_63; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_64 = io_sc2mac_wt_mask_64; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_65 = io_sc2mac_wt_mask_65; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_66 = io_sc2mac_wt_mask_66; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_67 = io_sc2mac_wt_mask_67; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_68 = io_sc2mac_wt_mask_68; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_69 = io_sc2mac_wt_mask_69; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_70 = io_sc2mac_wt_mask_70; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_71 = io_sc2mac_wt_mask_71; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_72 = io_sc2mac_wt_mask_72; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_73 = io_sc2mac_wt_mask_73; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_74 = io_sc2mac_wt_mask_74; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_75 = io_sc2mac_wt_mask_75; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_76 = io_sc2mac_wt_mask_76; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_77 = io_sc2mac_wt_mask_77; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_78 = io_sc2mac_wt_mask_78; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_79 = io_sc2mac_wt_mask_79; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_80 = io_sc2mac_wt_mask_80; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_81 = io_sc2mac_wt_mask_81; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_82 = io_sc2mac_wt_mask_82; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_83 = io_sc2mac_wt_mask_83; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_84 = io_sc2mac_wt_mask_84; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_85 = io_sc2mac_wt_mask_85; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_86 = io_sc2mac_wt_mask_86; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_87 = io_sc2mac_wt_mask_87; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_88 = io_sc2mac_wt_mask_88; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_89 = io_sc2mac_wt_mask_89; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_90 = io_sc2mac_wt_mask_90; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_91 = io_sc2mac_wt_mask_91; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_92 = io_sc2mac_wt_mask_92; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_93 = io_sc2mac_wt_mask_93; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_94 = io_sc2mac_wt_mask_94; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_95 = io_sc2mac_wt_mask_95; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_96 = io_sc2mac_wt_mask_96; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_97 = io_sc2mac_wt_mask_97; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_98 = io_sc2mac_wt_mask_98; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_99 = io_sc2mac_wt_mask_99; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_100 = io_sc2mac_wt_mask_100; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_101 = io_sc2mac_wt_mask_101; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_102 = io_sc2mac_wt_mask_102; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_103 = io_sc2mac_wt_mask_103; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_104 = io_sc2mac_wt_mask_104; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_105 = io_sc2mac_wt_mask_105; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_106 = io_sc2mac_wt_mask_106; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_107 = io_sc2mac_wt_mask_107; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_108 = io_sc2mac_wt_mask_108; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_109 = io_sc2mac_wt_mask_109; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_110 = io_sc2mac_wt_mask_110; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_111 = io_sc2mac_wt_mask_111; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_112 = io_sc2mac_wt_mask_112; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_113 = io_sc2mac_wt_mask_113; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_114 = io_sc2mac_wt_mask_114; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_115 = io_sc2mac_wt_mask_115; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_116 = io_sc2mac_wt_mask_116; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_117 = io_sc2mac_wt_mask_117; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_118 = io_sc2mac_wt_mask_118; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_119 = io_sc2mac_wt_mask_119; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_120 = io_sc2mac_wt_mask_120; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_121 = io_sc2mac_wt_mask_121; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_122 = io_sc2mac_wt_mask_122; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_123 = io_sc2mac_wt_mask_123; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_124 = io_sc2mac_wt_mask_124; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_125 = io_sc2mac_wt_mask_125; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_126 = io_sc2mac_wt_mask_126; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_mask_127 = io_sc2mac_wt_mask_127; // @[NV_NVDLA_CMAC_core.scala 60:31]
  assign u_rt_in_io_sc2mac_wt_sel_0 = io_sc2mac_wt_sel_0; // @[NV_NVDLA_CMAC_core.scala 62:30]
  assign u_rt_in_io_sc2mac_wt_pvld = io_sc2mac_wt_pvld; // @[NV_NVDLA_CMAC_core.scala 59:31]
  assign u_active_clock = clock;
  assign u_active_reset = reset;
  assign u_active_io_in_dat_data_0 = u_rt_in_io_in_dat_data_0; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_1 = u_rt_in_io_in_dat_data_1; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_2 = u_rt_in_io_in_dat_data_2; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_3 = u_rt_in_io_in_dat_data_3; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_4 = u_rt_in_io_in_dat_data_4; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_5 = u_rt_in_io_in_dat_data_5; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_6 = u_rt_in_io_in_dat_data_6; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_7 = u_rt_in_io_in_dat_data_7; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_8 = u_rt_in_io_in_dat_data_8; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_9 = u_rt_in_io_in_dat_data_9; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_10 = u_rt_in_io_in_dat_data_10; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_11 = u_rt_in_io_in_dat_data_11; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_12 = u_rt_in_io_in_dat_data_12; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_13 = u_rt_in_io_in_dat_data_13; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_14 = u_rt_in_io_in_dat_data_14; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_15 = u_rt_in_io_in_dat_data_15; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_16 = u_rt_in_io_in_dat_data_16; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_17 = u_rt_in_io_in_dat_data_17; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_18 = u_rt_in_io_in_dat_data_18; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_19 = u_rt_in_io_in_dat_data_19; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_20 = u_rt_in_io_in_dat_data_20; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_21 = u_rt_in_io_in_dat_data_21; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_22 = u_rt_in_io_in_dat_data_22; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_23 = u_rt_in_io_in_dat_data_23; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_24 = u_rt_in_io_in_dat_data_24; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_25 = u_rt_in_io_in_dat_data_25; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_26 = u_rt_in_io_in_dat_data_26; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_27 = u_rt_in_io_in_dat_data_27; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_28 = u_rt_in_io_in_dat_data_28; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_29 = u_rt_in_io_in_dat_data_29; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_30 = u_rt_in_io_in_dat_data_30; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_31 = u_rt_in_io_in_dat_data_31; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_32 = u_rt_in_io_in_dat_data_32; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_33 = u_rt_in_io_in_dat_data_33; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_34 = u_rt_in_io_in_dat_data_34; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_35 = u_rt_in_io_in_dat_data_35; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_36 = u_rt_in_io_in_dat_data_36; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_37 = u_rt_in_io_in_dat_data_37; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_38 = u_rt_in_io_in_dat_data_38; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_39 = u_rt_in_io_in_dat_data_39; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_40 = u_rt_in_io_in_dat_data_40; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_41 = u_rt_in_io_in_dat_data_41; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_42 = u_rt_in_io_in_dat_data_42; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_43 = u_rt_in_io_in_dat_data_43; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_44 = u_rt_in_io_in_dat_data_44; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_45 = u_rt_in_io_in_dat_data_45; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_46 = u_rt_in_io_in_dat_data_46; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_47 = u_rt_in_io_in_dat_data_47; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_48 = u_rt_in_io_in_dat_data_48; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_49 = u_rt_in_io_in_dat_data_49; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_50 = u_rt_in_io_in_dat_data_50; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_51 = u_rt_in_io_in_dat_data_51; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_52 = u_rt_in_io_in_dat_data_52; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_53 = u_rt_in_io_in_dat_data_53; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_54 = u_rt_in_io_in_dat_data_54; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_55 = u_rt_in_io_in_dat_data_55; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_56 = u_rt_in_io_in_dat_data_56; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_57 = u_rt_in_io_in_dat_data_57; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_58 = u_rt_in_io_in_dat_data_58; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_59 = u_rt_in_io_in_dat_data_59; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_60 = u_rt_in_io_in_dat_data_60; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_61 = u_rt_in_io_in_dat_data_61; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_62 = u_rt_in_io_in_dat_data_62; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_63 = u_rt_in_io_in_dat_data_63; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_64 = u_rt_in_io_in_dat_data_64; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_65 = u_rt_in_io_in_dat_data_65; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_66 = u_rt_in_io_in_dat_data_66; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_67 = u_rt_in_io_in_dat_data_67; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_68 = u_rt_in_io_in_dat_data_68; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_69 = u_rt_in_io_in_dat_data_69; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_70 = u_rt_in_io_in_dat_data_70; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_71 = u_rt_in_io_in_dat_data_71; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_72 = u_rt_in_io_in_dat_data_72; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_73 = u_rt_in_io_in_dat_data_73; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_74 = u_rt_in_io_in_dat_data_74; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_75 = u_rt_in_io_in_dat_data_75; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_76 = u_rt_in_io_in_dat_data_76; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_77 = u_rt_in_io_in_dat_data_77; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_78 = u_rt_in_io_in_dat_data_78; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_79 = u_rt_in_io_in_dat_data_79; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_80 = u_rt_in_io_in_dat_data_80; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_81 = u_rt_in_io_in_dat_data_81; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_82 = u_rt_in_io_in_dat_data_82; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_83 = u_rt_in_io_in_dat_data_83; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_84 = u_rt_in_io_in_dat_data_84; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_85 = u_rt_in_io_in_dat_data_85; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_86 = u_rt_in_io_in_dat_data_86; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_87 = u_rt_in_io_in_dat_data_87; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_88 = u_rt_in_io_in_dat_data_88; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_89 = u_rt_in_io_in_dat_data_89; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_90 = u_rt_in_io_in_dat_data_90; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_91 = u_rt_in_io_in_dat_data_91; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_92 = u_rt_in_io_in_dat_data_92; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_93 = u_rt_in_io_in_dat_data_93; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_94 = u_rt_in_io_in_dat_data_94; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_95 = u_rt_in_io_in_dat_data_95; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_96 = u_rt_in_io_in_dat_data_96; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_97 = u_rt_in_io_in_dat_data_97; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_98 = u_rt_in_io_in_dat_data_98; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_99 = u_rt_in_io_in_dat_data_99; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_100 = u_rt_in_io_in_dat_data_100; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_101 = u_rt_in_io_in_dat_data_101; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_102 = u_rt_in_io_in_dat_data_102; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_103 = u_rt_in_io_in_dat_data_103; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_104 = u_rt_in_io_in_dat_data_104; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_105 = u_rt_in_io_in_dat_data_105; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_106 = u_rt_in_io_in_dat_data_106; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_107 = u_rt_in_io_in_dat_data_107; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_108 = u_rt_in_io_in_dat_data_108; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_109 = u_rt_in_io_in_dat_data_109; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_110 = u_rt_in_io_in_dat_data_110; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_111 = u_rt_in_io_in_dat_data_111; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_112 = u_rt_in_io_in_dat_data_112; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_113 = u_rt_in_io_in_dat_data_113; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_114 = u_rt_in_io_in_dat_data_114; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_115 = u_rt_in_io_in_dat_data_115; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_116 = u_rt_in_io_in_dat_data_116; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_117 = u_rt_in_io_in_dat_data_117; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_118 = u_rt_in_io_in_dat_data_118; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_119 = u_rt_in_io_in_dat_data_119; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_120 = u_rt_in_io_in_dat_data_120; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_121 = u_rt_in_io_in_dat_data_121; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_122 = u_rt_in_io_in_dat_data_122; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_123 = u_rt_in_io_in_dat_data_123; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_124 = u_rt_in_io_in_dat_data_124; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_125 = u_rt_in_io_in_dat_data_125; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_126 = u_rt_in_io_in_dat_data_126; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_data_127 = u_rt_in_io_in_dat_data_127; // @[NV_NVDLA_CMAC_core.scala 86:29]
  assign u_active_io_in_dat_mask_0 = u_rt_in_io_in_dat_mask_0; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_1 = u_rt_in_io_in_dat_mask_1; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_2 = u_rt_in_io_in_dat_mask_2; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_3 = u_rt_in_io_in_dat_mask_3; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_4 = u_rt_in_io_in_dat_mask_4; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_5 = u_rt_in_io_in_dat_mask_5; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_6 = u_rt_in_io_in_dat_mask_6; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_7 = u_rt_in_io_in_dat_mask_7; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_8 = u_rt_in_io_in_dat_mask_8; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_9 = u_rt_in_io_in_dat_mask_9; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_10 = u_rt_in_io_in_dat_mask_10; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_11 = u_rt_in_io_in_dat_mask_11; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_12 = u_rt_in_io_in_dat_mask_12; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_13 = u_rt_in_io_in_dat_mask_13; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_14 = u_rt_in_io_in_dat_mask_14; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_15 = u_rt_in_io_in_dat_mask_15; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_16 = u_rt_in_io_in_dat_mask_16; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_17 = u_rt_in_io_in_dat_mask_17; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_18 = u_rt_in_io_in_dat_mask_18; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_19 = u_rt_in_io_in_dat_mask_19; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_20 = u_rt_in_io_in_dat_mask_20; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_21 = u_rt_in_io_in_dat_mask_21; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_22 = u_rt_in_io_in_dat_mask_22; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_23 = u_rt_in_io_in_dat_mask_23; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_24 = u_rt_in_io_in_dat_mask_24; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_25 = u_rt_in_io_in_dat_mask_25; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_26 = u_rt_in_io_in_dat_mask_26; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_27 = u_rt_in_io_in_dat_mask_27; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_28 = u_rt_in_io_in_dat_mask_28; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_29 = u_rt_in_io_in_dat_mask_29; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_30 = u_rt_in_io_in_dat_mask_30; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_31 = u_rt_in_io_in_dat_mask_31; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_32 = u_rt_in_io_in_dat_mask_32; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_33 = u_rt_in_io_in_dat_mask_33; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_34 = u_rt_in_io_in_dat_mask_34; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_35 = u_rt_in_io_in_dat_mask_35; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_36 = u_rt_in_io_in_dat_mask_36; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_37 = u_rt_in_io_in_dat_mask_37; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_38 = u_rt_in_io_in_dat_mask_38; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_39 = u_rt_in_io_in_dat_mask_39; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_40 = u_rt_in_io_in_dat_mask_40; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_41 = u_rt_in_io_in_dat_mask_41; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_42 = u_rt_in_io_in_dat_mask_42; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_43 = u_rt_in_io_in_dat_mask_43; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_44 = u_rt_in_io_in_dat_mask_44; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_45 = u_rt_in_io_in_dat_mask_45; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_46 = u_rt_in_io_in_dat_mask_46; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_47 = u_rt_in_io_in_dat_mask_47; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_48 = u_rt_in_io_in_dat_mask_48; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_49 = u_rt_in_io_in_dat_mask_49; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_50 = u_rt_in_io_in_dat_mask_50; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_51 = u_rt_in_io_in_dat_mask_51; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_52 = u_rt_in_io_in_dat_mask_52; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_53 = u_rt_in_io_in_dat_mask_53; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_54 = u_rt_in_io_in_dat_mask_54; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_55 = u_rt_in_io_in_dat_mask_55; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_56 = u_rt_in_io_in_dat_mask_56; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_57 = u_rt_in_io_in_dat_mask_57; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_58 = u_rt_in_io_in_dat_mask_58; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_59 = u_rt_in_io_in_dat_mask_59; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_60 = u_rt_in_io_in_dat_mask_60; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_61 = u_rt_in_io_in_dat_mask_61; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_62 = u_rt_in_io_in_dat_mask_62; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_63 = u_rt_in_io_in_dat_mask_63; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_64 = u_rt_in_io_in_dat_mask_64; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_65 = u_rt_in_io_in_dat_mask_65; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_66 = u_rt_in_io_in_dat_mask_66; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_67 = u_rt_in_io_in_dat_mask_67; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_68 = u_rt_in_io_in_dat_mask_68; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_69 = u_rt_in_io_in_dat_mask_69; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_70 = u_rt_in_io_in_dat_mask_70; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_71 = u_rt_in_io_in_dat_mask_71; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_72 = u_rt_in_io_in_dat_mask_72; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_73 = u_rt_in_io_in_dat_mask_73; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_74 = u_rt_in_io_in_dat_mask_74; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_75 = u_rt_in_io_in_dat_mask_75; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_76 = u_rt_in_io_in_dat_mask_76; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_77 = u_rt_in_io_in_dat_mask_77; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_78 = u_rt_in_io_in_dat_mask_78; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_79 = u_rt_in_io_in_dat_mask_79; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_80 = u_rt_in_io_in_dat_mask_80; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_81 = u_rt_in_io_in_dat_mask_81; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_82 = u_rt_in_io_in_dat_mask_82; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_83 = u_rt_in_io_in_dat_mask_83; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_84 = u_rt_in_io_in_dat_mask_84; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_85 = u_rt_in_io_in_dat_mask_85; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_86 = u_rt_in_io_in_dat_mask_86; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_87 = u_rt_in_io_in_dat_mask_87; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_88 = u_rt_in_io_in_dat_mask_88; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_89 = u_rt_in_io_in_dat_mask_89; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_90 = u_rt_in_io_in_dat_mask_90; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_91 = u_rt_in_io_in_dat_mask_91; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_92 = u_rt_in_io_in_dat_mask_92; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_93 = u_rt_in_io_in_dat_mask_93; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_94 = u_rt_in_io_in_dat_mask_94; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_95 = u_rt_in_io_in_dat_mask_95; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_96 = u_rt_in_io_in_dat_mask_96; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_97 = u_rt_in_io_in_dat_mask_97; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_98 = u_rt_in_io_in_dat_mask_98; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_99 = u_rt_in_io_in_dat_mask_99; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_100 = u_rt_in_io_in_dat_mask_100; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_101 = u_rt_in_io_in_dat_mask_101; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_102 = u_rt_in_io_in_dat_mask_102; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_103 = u_rt_in_io_in_dat_mask_103; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_104 = u_rt_in_io_in_dat_mask_104; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_105 = u_rt_in_io_in_dat_mask_105; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_106 = u_rt_in_io_in_dat_mask_106; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_107 = u_rt_in_io_in_dat_mask_107; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_108 = u_rt_in_io_in_dat_mask_108; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_109 = u_rt_in_io_in_dat_mask_109; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_110 = u_rt_in_io_in_dat_mask_110; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_111 = u_rt_in_io_in_dat_mask_111; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_112 = u_rt_in_io_in_dat_mask_112; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_113 = u_rt_in_io_in_dat_mask_113; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_114 = u_rt_in_io_in_dat_mask_114; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_115 = u_rt_in_io_in_dat_mask_115; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_116 = u_rt_in_io_in_dat_mask_116; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_117 = u_rt_in_io_in_dat_mask_117; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_118 = u_rt_in_io_in_dat_mask_118; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_119 = u_rt_in_io_in_dat_mask_119; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_120 = u_rt_in_io_in_dat_mask_120; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_121 = u_rt_in_io_in_dat_mask_121; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_122 = u_rt_in_io_in_dat_mask_122; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_123 = u_rt_in_io_in_dat_mask_123; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_124 = u_rt_in_io_in_dat_mask_124; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_125 = u_rt_in_io_in_dat_mask_125; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_126 = u_rt_in_io_in_dat_mask_126; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_mask_127 = u_rt_in_io_in_dat_mask_127; // @[NV_NVDLA_CMAC_core.scala 85:29]
  assign u_active_io_in_dat_pvld = u_rt_in_io_in_dat_pvld; // @[NV_NVDLA_CMAC_core.scala 84:29]
  assign u_active_io_in_dat_stripe_st = u_rt_in_io_in_dat_stripe_st; // @[NV_NVDLA_CMAC_core.scala 88:34]
  assign u_active_io_in_dat_stripe_end = u_rt_in_io_in_dat_stripe_end; // @[NV_NVDLA_CMAC_core.scala 87:35]
  assign u_active_io_in_wt_data_0 = u_rt_in_io_in_wt_data_0; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_1 = u_rt_in_io_in_wt_data_1; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_2 = u_rt_in_io_in_wt_data_2; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_3 = u_rt_in_io_in_wt_data_3; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_4 = u_rt_in_io_in_wt_data_4; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_5 = u_rt_in_io_in_wt_data_5; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_6 = u_rt_in_io_in_wt_data_6; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_7 = u_rt_in_io_in_wt_data_7; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_8 = u_rt_in_io_in_wt_data_8; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_9 = u_rt_in_io_in_wt_data_9; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_10 = u_rt_in_io_in_wt_data_10; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_11 = u_rt_in_io_in_wt_data_11; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_12 = u_rt_in_io_in_wt_data_12; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_13 = u_rt_in_io_in_wt_data_13; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_14 = u_rt_in_io_in_wt_data_14; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_15 = u_rt_in_io_in_wt_data_15; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_16 = u_rt_in_io_in_wt_data_16; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_17 = u_rt_in_io_in_wt_data_17; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_18 = u_rt_in_io_in_wt_data_18; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_19 = u_rt_in_io_in_wt_data_19; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_20 = u_rt_in_io_in_wt_data_20; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_21 = u_rt_in_io_in_wt_data_21; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_22 = u_rt_in_io_in_wt_data_22; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_23 = u_rt_in_io_in_wt_data_23; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_24 = u_rt_in_io_in_wt_data_24; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_25 = u_rt_in_io_in_wt_data_25; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_26 = u_rt_in_io_in_wt_data_26; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_27 = u_rt_in_io_in_wt_data_27; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_28 = u_rt_in_io_in_wt_data_28; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_29 = u_rt_in_io_in_wt_data_29; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_30 = u_rt_in_io_in_wt_data_30; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_31 = u_rt_in_io_in_wt_data_31; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_32 = u_rt_in_io_in_wt_data_32; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_33 = u_rt_in_io_in_wt_data_33; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_34 = u_rt_in_io_in_wt_data_34; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_35 = u_rt_in_io_in_wt_data_35; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_36 = u_rt_in_io_in_wt_data_36; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_37 = u_rt_in_io_in_wt_data_37; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_38 = u_rt_in_io_in_wt_data_38; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_39 = u_rt_in_io_in_wt_data_39; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_40 = u_rt_in_io_in_wt_data_40; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_41 = u_rt_in_io_in_wt_data_41; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_42 = u_rt_in_io_in_wt_data_42; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_43 = u_rt_in_io_in_wt_data_43; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_44 = u_rt_in_io_in_wt_data_44; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_45 = u_rt_in_io_in_wt_data_45; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_46 = u_rt_in_io_in_wt_data_46; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_47 = u_rt_in_io_in_wt_data_47; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_48 = u_rt_in_io_in_wt_data_48; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_49 = u_rt_in_io_in_wt_data_49; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_50 = u_rt_in_io_in_wt_data_50; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_51 = u_rt_in_io_in_wt_data_51; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_52 = u_rt_in_io_in_wt_data_52; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_53 = u_rt_in_io_in_wt_data_53; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_54 = u_rt_in_io_in_wt_data_54; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_55 = u_rt_in_io_in_wt_data_55; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_56 = u_rt_in_io_in_wt_data_56; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_57 = u_rt_in_io_in_wt_data_57; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_58 = u_rt_in_io_in_wt_data_58; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_59 = u_rt_in_io_in_wt_data_59; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_60 = u_rt_in_io_in_wt_data_60; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_61 = u_rt_in_io_in_wt_data_61; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_62 = u_rt_in_io_in_wt_data_62; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_63 = u_rt_in_io_in_wt_data_63; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_64 = u_rt_in_io_in_wt_data_64; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_65 = u_rt_in_io_in_wt_data_65; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_66 = u_rt_in_io_in_wt_data_66; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_67 = u_rt_in_io_in_wt_data_67; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_68 = u_rt_in_io_in_wt_data_68; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_69 = u_rt_in_io_in_wt_data_69; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_70 = u_rt_in_io_in_wt_data_70; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_71 = u_rt_in_io_in_wt_data_71; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_72 = u_rt_in_io_in_wt_data_72; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_73 = u_rt_in_io_in_wt_data_73; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_74 = u_rt_in_io_in_wt_data_74; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_75 = u_rt_in_io_in_wt_data_75; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_76 = u_rt_in_io_in_wt_data_76; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_77 = u_rt_in_io_in_wt_data_77; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_78 = u_rt_in_io_in_wt_data_78; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_79 = u_rt_in_io_in_wt_data_79; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_80 = u_rt_in_io_in_wt_data_80; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_81 = u_rt_in_io_in_wt_data_81; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_82 = u_rt_in_io_in_wt_data_82; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_83 = u_rt_in_io_in_wt_data_83; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_84 = u_rt_in_io_in_wt_data_84; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_85 = u_rt_in_io_in_wt_data_85; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_86 = u_rt_in_io_in_wt_data_86; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_87 = u_rt_in_io_in_wt_data_87; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_88 = u_rt_in_io_in_wt_data_88; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_89 = u_rt_in_io_in_wt_data_89; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_90 = u_rt_in_io_in_wt_data_90; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_91 = u_rt_in_io_in_wt_data_91; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_92 = u_rt_in_io_in_wt_data_92; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_93 = u_rt_in_io_in_wt_data_93; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_94 = u_rt_in_io_in_wt_data_94; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_95 = u_rt_in_io_in_wt_data_95; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_96 = u_rt_in_io_in_wt_data_96; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_97 = u_rt_in_io_in_wt_data_97; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_98 = u_rt_in_io_in_wt_data_98; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_99 = u_rt_in_io_in_wt_data_99; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_100 = u_rt_in_io_in_wt_data_100; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_101 = u_rt_in_io_in_wt_data_101; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_102 = u_rt_in_io_in_wt_data_102; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_103 = u_rt_in_io_in_wt_data_103; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_104 = u_rt_in_io_in_wt_data_104; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_105 = u_rt_in_io_in_wt_data_105; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_106 = u_rt_in_io_in_wt_data_106; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_107 = u_rt_in_io_in_wt_data_107; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_108 = u_rt_in_io_in_wt_data_108; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_109 = u_rt_in_io_in_wt_data_109; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_110 = u_rt_in_io_in_wt_data_110; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_111 = u_rt_in_io_in_wt_data_111; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_112 = u_rt_in_io_in_wt_data_112; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_113 = u_rt_in_io_in_wt_data_113; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_114 = u_rt_in_io_in_wt_data_114; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_115 = u_rt_in_io_in_wt_data_115; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_116 = u_rt_in_io_in_wt_data_116; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_117 = u_rt_in_io_in_wt_data_117; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_118 = u_rt_in_io_in_wt_data_118; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_119 = u_rt_in_io_in_wt_data_119; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_120 = u_rt_in_io_in_wt_data_120; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_121 = u_rt_in_io_in_wt_data_121; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_122 = u_rt_in_io_in_wt_data_122; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_123 = u_rt_in_io_in_wt_data_123; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_124 = u_rt_in_io_in_wt_data_124; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_125 = u_rt_in_io_in_wt_data_125; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_126 = u_rt_in_io_in_wt_data_126; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_data_127 = u_rt_in_io_in_wt_data_127; // @[NV_NVDLA_CMAC_core.scala 92:28]
  assign u_active_io_in_wt_mask_0 = u_rt_in_io_in_wt_mask_0; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_1 = u_rt_in_io_in_wt_mask_1; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_2 = u_rt_in_io_in_wt_mask_2; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_3 = u_rt_in_io_in_wt_mask_3; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_4 = u_rt_in_io_in_wt_mask_4; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_5 = u_rt_in_io_in_wt_mask_5; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_6 = u_rt_in_io_in_wt_mask_6; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_7 = u_rt_in_io_in_wt_mask_7; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_8 = u_rt_in_io_in_wt_mask_8; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_9 = u_rt_in_io_in_wt_mask_9; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_10 = u_rt_in_io_in_wt_mask_10; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_11 = u_rt_in_io_in_wt_mask_11; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_12 = u_rt_in_io_in_wt_mask_12; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_13 = u_rt_in_io_in_wt_mask_13; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_14 = u_rt_in_io_in_wt_mask_14; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_15 = u_rt_in_io_in_wt_mask_15; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_16 = u_rt_in_io_in_wt_mask_16; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_17 = u_rt_in_io_in_wt_mask_17; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_18 = u_rt_in_io_in_wt_mask_18; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_19 = u_rt_in_io_in_wt_mask_19; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_20 = u_rt_in_io_in_wt_mask_20; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_21 = u_rt_in_io_in_wt_mask_21; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_22 = u_rt_in_io_in_wt_mask_22; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_23 = u_rt_in_io_in_wt_mask_23; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_24 = u_rt_in_io_in_wt_mask_24; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_25 = u_rt_in_io_in_wt_mask_25; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_26 = u_rt_in_io_in_wt_mask_26; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_27 = u_rt_in_io_in_wt_mask_27; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_28 = u_rt_in_io_in_wt_mask_28; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_29 = u_rt_in_io_in_wt_mask_29; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_30 = u_rt_in_io_in_wt_mask_30; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_31 = u_rt_in_io_in_wt_mask_31; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_32 = u_rt_in_io_in_wt_mask_32; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_33 = u_rt_in_io_in_wt_mask_33; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_34 = u_rt_in_io_in_wt_mask_34; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_35 = u_rt_in_io_in_wt_mask_35; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_36 = u_rt_in_io_in_wt_mask_36; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_37 = u_rt_in_io_in_wt_mask_37; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_38 = u_rt_in_io_in_wt_mask_38; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_39 = u_rt_in_io_in_wt_mask_39; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_40 = u_rt_in_io_in_wt_mask_40; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_41 = u_rt_in_io_in_wt_mask_41; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_42 = u_rt_in_io_in_wt_mask_42; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_43 = u_rt_in_io_in_wt_mask_43; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_44 = u_rt_in_io_in_wt_mask_44; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_45 = u_rt_in_io_in_wt_mask_45; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_46 = u_rt_in_io_in_wt_mask_46; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_47 = u_rt_in_io_in_wt_mask_47; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_48 = u_rt_in_io_in_wt_mask_48; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_49 = u_rt_in_io_in_wt_mask_49; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_50 = u_rt_in_io_in_wt_mask_50; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_51 = u_rt_in_io_in_wt_mask_51; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_52 = u_rt_in_io_in_wt_mask_52; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_53 = u_rt_in_io_in_wt_mask_53; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_54 = u_rt_in_io_in_wt_mask_54; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_55 = u_rt_in_io_in_wt_mask_55; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_56 = u_rt_in_io_in_wt_mask_56; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_57 = u_rt_in_io_in_wt_mask_57; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_58 = u_rt_in_io_in_wt_mask_58; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_59 = u_rt_in_io_in_wt_mask_59; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_60 = u_rt_in_io_in_wt_mask_60; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_61 = u_rt_in_io_in_wt_mask_61; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_62 = u_rt_in_io_in_wt_mask_62; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_63 = u_rt_in_io_in_wt_mask_63; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_64 = u_rt_in_io_in_wt_mask_64; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_65 = u_rt_in_io_in_wt_mask_65; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_66 = u_rt_in_io_in_wt_mask_66; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_67 = u_rt_in_io_in_wt_mask_67; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_68 = u_rt_in_io_in_wt_mask_68; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_69 = u_rt_in_io_in_wt_mask_69; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_70 = u_rt_in_io_in_wt_mask_70; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_71 = u_rt_in_io_in_wt_mask_71; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_72 = u_rt_in_io_in_wt_mask_72; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_73 = u_rt_in_io_in_wt_mask_73; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_74 = u_rt_in_io_in_wt_mask_74; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_75 = u_rt_in_io_in_wt_mask_75; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_76 = u_rt_in_io_in_wt_mask_76; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_77 = u_rt_in_io_in_wt_mask_77; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_78 = u_rt_in_io_in_wt_mask_78; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_79 = u_rt_in_io_in_wt_mask_79; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_80 = u_rt_in_io_in_wt_mask_80; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_81 = u_rt_in_io_in_wt_mask_81; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_82 = u_rt_in_io_in_wt_mask_82; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_83 = u_rt_in_io_in_wt_mask_83; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_84 = u_rt_in_io_in_wt_mask_84; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_85 = u_rt_in_io_in_wt_mask_85; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_86 = u_rt_in_io_in_wt_mask_86; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_87 = u_rt_in_io_in_wt_mask_87; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_88 = u_rt_in_io_in_wt_mask_88; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_89 = u_rt_in_io_in_wt_mask_89; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_90 = u_rt_in_io_in_wt_mask_90; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_91 = u_rt_in_io_in_wt_mask_91; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_92 = u_rt_in_io_in_wt_mask_92; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_93 = u_rt_in_io_in_wt_mask_93; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_94 = u_rt_in_io_in_wt_mask_94; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_95 = u_rt_in_io_in_wt_mask_95; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_96 = u_rt_in_io_in_wt_mask_96; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_97 = u_rt_in_io_in_wt_mask_97; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_98 = u_rt_in_io_in_wt_mask_98; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_99 = u_rt_in_io_in_wt_mask_99; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_100 = u_rt_in_io_in_wt_mask_100; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_101 = u_rt_in_io_in_wt_mask_101; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_102 = u_rt_in_io_in_wt_mask_102; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_103 = u_rt_in_io_in_wt_mask_103; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_104 = u_rt_in_io_in_wt_mask_104; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_105 = u_rt_in_io_in_wt_mask_105; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_106 = u_rt_in_io_in_wt_mask_106; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_107 = u_rt_in_io_in_wt_mask_107; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_108 = u_rt_in_io_in_wt_mask_108; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_109 = u_rt_in_io_in_wt_mask_109; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_110 = u_rt_in_io_in_wt_mask_110; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_111 = u_rt_in_io_in_wt_mask_111; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_112 = u_rt_in_io_in_wt_mask_112; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_113 = u_rt_in_io_in_wt_mask_113; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_114 = u_rt_in_io_in_wt_mask_114; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_115 = u_rt_in_io_in_wt_mask_115; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_116 = u_rt_in_io_in_wt_mask_116; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_117 = u_rt_in_io_in_wt_mask_117; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_118 = u_rt_in_io_in_wt_mask_118; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_119 = u_rt_in_io_in_wt_mask_119; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_120 = u_rt_in_io_in_wt_mask_120; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_121 = u_rt_in_io_in_wt_mask_121; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_122 = u_rt_in_io_in_wt_mask_122; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_123 = u_rt_in_io_in_wt_mask_123; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_124 = u_rt_in_io_in_wt_mask_124; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_125 = u_rt_in_io_in_wt_mask_125; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_126 = u_rt_in_io_in_wt_mask_126; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_mask_127 = u_rt_in_io_in_wt_mask_127; // @[NV_NVDLA_CMAC_core.scala 91:28]
  assign u_active_io_in_wt_pvld = u_rt_in_io_in_wt_pvld; // @[NV_NVDLA_CMAC_core.scala 90:28]
  assign u_active_io_in_wt_sel_0 = u_rt_in_io_in_wt_sel_0; // @[NV_NVDLA_CMAC_core.scala 93:27]
  assign NV_NVDLA_CMAC_CORE_mac_clock = clock;
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_0 = u_active_io_dat_actv_data_0_0; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_1 = u_active_io_dat_actv_data_0_1; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_2 = u_active_io_dat_actv_data_0_2; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_3 = u_active_io_dat_actv_data_0_3; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_4 = u_active_io_dat_actv_data_0_4; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_5 = u_active_io_dat_actv_data_0_5; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_6 = u_active_io_dat_actv_data_0_6; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_7 = u_active_io_dat_actv_data_0_7; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_8 = u_active_io_dat_actv_data_0_8; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_9 = u_active_io_dat_actv_data_0_9; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_10 = u_active_io_dat_actv_data_0_10; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_11 = u_active_io_dat_actv_data_0_11; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_12 = u_active_io_dat_actv_data_0_12; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_13 = u_active_io_dat_actv_data_0_13; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_14 = u_active_io_dat_actv_data_0_14; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_15 = u_active_io_dat_actv_data_0_15; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_16 = u_active_io_dat_actv_data_0_16; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_17 = u_active_io_dat_actv_data_0_17; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_18 = u_active_io_dat_actv_data_0_18; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_19 = u_active_io_dat_actv_data_0_19; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_20 = u_active_io_dat_actv_data_0_20; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_21 = u_active_io_dat_actv_data_0_21; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_22 = u_active_io_dat_actv_data_0_22; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_23 = u_active_io_dat_actv_data_0_23; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_24 = u_active_io_dat_actv_data_0_24; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_25 = u_active_io_dat_actv_data_0_25; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_26 = u_active_io_dat_actv_data_0_26; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_27 = u_active_io_dat_actv_data_0_27; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_28 = u_active_io_dat_actv_data_0_28; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_29 = u_active_io_dat_actv_data_0_29; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_30 = u_active_io_dat_actv_data_0_30; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_31 = u_active_io_dat_actv_data_0_31; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_32 = u_active_io_dat_actv_data_0_32; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_33 = u_active_io_dat_actv_data_0_33; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_34 = u_active_io_dat_actv_data_0_34; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_35 = u_active_io_dat_actv_data_0_35; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_36 = u_active_io_dat_actv_data_0_36; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_37 = u_active_io_dat_actv_data_0_37; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_38 = u_active_io_dat_actv_data_0_38; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_39 = u_active_io_dat_actv_data_0_39; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_40 = u_active_io_dat_actv_data_0_40; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_41 = u_active_io_dat_actv_data_0_41; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_42 = u_active_io_dat_actv_data_0_42; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_43 = u_active_io_dat_actv_data_0_43; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_44 = u_active_io_dat_actv_data_0_44; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_45 = u_active_io_dat_actv_data_0_45; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_46 = u_active_io_dat_actv_data_0_46; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_47 = u_active_io_dat_actv_data_0_47; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_48 = u_active_io_dat_actv_data_0_48; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_49 = u_active_io_dat_actv_data_0_49; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_50 = u_active_io_dat_actv_data_0_50; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_51 = u_active_io_dat_actv_data_0_51; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_52 = u_active_io_dat_actv_data_0_52; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_53 = u_active_io_dat_actv_data_0_53; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_54 = u_active_io_dat_actv_data_0_54; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_55 = u_active_io_dat_actv_data_0_55; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_56 = u_active_io_dat_actv_data_0_56; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_57 = u_active_io_dat_actv_data_0_57; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_58 = u_active_io_dat_actv_data_0_58; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_59 = u_active_io_dat_actv_data_0_59; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_60 = u_active_io_dat_actv_data_0_60; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_61 = u_active_io_dat_actv_data_0_61; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_62 = u_active_io_dat_actv_data_0_62; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_63 = u_active_io_dat_actv_data_0_63; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_64 = u_active_io_dat_actv_data_0_64; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_65 = u_active_io_dat_actv_data_0_65; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_66 = u_active_io_dat_actv_data_0_66; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_67 = u_active_io_dat_actv_data_0_67; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_68 = u_active_io_dat_actv_data_0_68; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_69 = u_active_io_dat_actv_data_0_69; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_70 = u_active_io_dat_actv_data_0_70; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_71 = u_active_io_dat_actv_data_0_71; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_72 = u_active_io_dat_actv_data_0_72; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_73 = u_active_io_dat_actv_data_0_73; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_74 = u_active_io_dat_actv_data_0_74; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_75 = u_active_io_dat_actv_data_0_75; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_76 = u_active_io_dat_actv_data_0_76; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_77 = u_active_io_dat_actv_data_0_77; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_78 = u_active_io_dat_actv_data_0_78; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_79 = u_active_io_dat_actv_data_0_79; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_80 = u_active_io_dat_actv_data_0_80; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_81 = u_active_io_dat_actv_data_0_81; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_82 = u_active_io_dat_actv_data_0_82; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_83 = u_active_io_dat_actv_data_0_83; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_84 = u_active_io_dat_actv_data_0_84; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_85 = u_active_io_dat_actv_data_0_85; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_86 = u_active_io_dat_actv_data_0_86; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_87 = u_active_io_dat_actv_data_0_87; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_88 = u_active_io_dat_actv_data_0_88; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_89 = u_active_io_dat_actv_data_0_89; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_90 = u_active_io_dat_actv_data_0_90; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_91 = u_active_io_dat_actv_data_0_91; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_92 = u_active_io_dat_actv_data_0_92; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_93 = u_active_io_dat_actv_data_0_93; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_94 = u_active_io_dat_actv_data_0_94; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_95 = u_active_io_dat_actv_data_0_95; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_96 = u_active_io_dat_actv_data_0_96; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_97 = u_active_io_dat_actv_data_0_97; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_98 = u_active_io_dat_actv_data_0_98; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_99 = u_active_io_dat_actv_data_0_99; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_100 = u_active_io_dat_actv_data_0_100; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_101 = u_active_io_dat_actv_data_0_101; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_102 = u_active_io_dat_actv_data_0_102; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_103 = u_active_io_dat_actv_data_0_103; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_104 = u_active_io_dat_actv_data_0_104; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_105 = u_active_io_dat_actv_data_0_105; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_106 = u_active_io_dat_actv_data_0_106; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_107 = u_active_io_dat_actv_data_0_107; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_108 = u_active_io_dat_actv_data_0_108; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_109 = u_active_io_dat_actv_data_0_109; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_110 = u_active_io_dat_actv_data_0_110; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_111 = u_active_io_dat_actv_data_0_111; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_112 = u_active_io_dat_actv_data_0_112; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_113 = u_active_io_dat_actv_data_0_113; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_114 = u_active_io_dat_actv_data_0_114; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_115 = u_active_io_dat_actv_data_0_115; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_116 = u_active_io_dat_actv_data_0_116; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_117 = u_active_io_dat_actv_data_0_117; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_118 = u_active_io_dat_actv_data_0_118; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_119 = u_active_io_dat_actv_data_0_119; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_120 = u_active_io_dat_actv_data_0_120; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_121 = u_active_io_dat_actv_data_0_121; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_122 = u_active_io_dat_actv_data_0_122; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_123 = u_active_io_dat_actv_data_0_123; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_124 = u_active_io_dat_actv_data_0_124; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_125 = u_active_io_dat_actv_data_0_125; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_126 = u_active_io_dat_actv_data_0_126; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_data_127 = u_active_io_dat_actv_data_0_127; // @[NV_NVDLA_CMAC_core.scala 116:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_0 = u_active_io_dat_actv_nz_0_0; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_1 = u_active_io_dat_actv_nz_0_1; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_2 = u_active_io_dat_actv_nz_0_2; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_3 = u_active_io_dat_actv_nz_0_3; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_4 = u_active_io_dat_actv_nz_0_4; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_5 = u_active_io_dat_actv_nz_0_5; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_6 = u_active_io_dat_actv_nz_0_6; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_7 = u_active_io_dat_actv_nz_0_7; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_8 = u_active_io_dat_actv_nz_0_8; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_9 = u_active_io_dat_actv_nz_0_9; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_10 = u_active_io_dat_actv_nz_0_10; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_11 = u_active_io_dat_actv_nz_0_11; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_12 = u_active_io_dat_actv_nz_0_12; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_13 = u_active_io_dat_actv_nz_0_13; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_14 = u_active_io_dat_actv_nz_0_14; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_15 = u_active_io_dat_actv_nz_0_15; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_16 = u_active_io_dat_actv_nz_0_16; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_17 = u_active_io_dat_actv_nz_0_17; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_18 = u_active_io_dat_actv_nz_0_18; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_19 = u_active_io_dat_actv_nz_0_19; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_20 = u_active_io_dat_actv_nz_0_20; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_21 = u_active_io_dat_actv_nz_0_21; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_22 = u_active_io_dat_actv_nz_0_22; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_23 = u_active_io_dat_actv_nz_0_23; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_24 = u_active_io_dat_actv_nz_0_24; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_25 = u_active_io_dat_actv_nz_0_25; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_26 = u_active_io_dat_actv_nz_0_26; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_27 = u_active_io_dat_actv_nz_0_27; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_28 = u_active_io_dat_actv_nz_0_28; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_29 = u_active_io_dat_actv_nz_0_29; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_30 = u_active_io_dat_actv_nz_0_30; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_31 = u_active_io_dat_actv_nz_0_31; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_32 = u_active_io_dat_actv_nz_0_32; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_33 = u_active_io_dat_actv_nz_0_33; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_34 = u_active_io_dat_actv_nz_0_34; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_35 = u_active_io_dat_actv_nz_0_35; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_36 = u_active_io_dat_actv_nz_0_36; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_37 = u_active_io_dat_actv_nz_0_37; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_38 = u_active_io_dat_actv_nz_0_38; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_39 = u_active_io_dat_actv_nz_0_39; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_40 = u_active_io_dat_actv_nz_0_40; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_41 = u_active_io_dat_actv_nz_0_41; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_42 = u_active_io_dat_actv_nz_0_42; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_43 = u_active_io_dat_actv_nz_0_43; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_44 = u_active_io_dat_actv_nz_0_44; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_45 = u_active_io_dat_actv_nz_0_45; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_46 = u_active_io_dat_actv_nz_0_46; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_47 = u_active_io_dat_actv_nz_0_47; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_48 = u_active_io_dat_actv_nz_0_48; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_49 = u_active_io_dat_actv_nz_0_49; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_50 = u_active_io_dat_actv_nz_0_50; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_51 = u_active_io_dat_actv_nz_0_51; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_52 = u_active_io_dat_actv_nz_0_52; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_53 = u_active_io_dat_actv_nz_0_53; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_54 = u_active_io_dat_actv_nz_0_54; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_55 = u_active_io_dat_actv_nz_0_55; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_56 = u_active_io_dat_actv_nz_0_56; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_57 = u_active_io_dat_actv_nz_0_57; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_58 = u_active_io_dat_actv_nz_0_58; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_59 = u_active_io_dat_actv_nz_0_59; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_60 = u_active_io_dat_actv_nz_0_60; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_61 = u_active_io_dat_actv_nz_0_61; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_62 = u_active_io_dat_actv_nz_0_62; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_63 = u_active_io_dat_actv_nz_0_63; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_64 = u_active_io_dat_actv_nz_0_64; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_65 = u_active_io_dat_actv_nz_0_65; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_66 = u_active_io_dat_actv_nz_0_66; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_67 = u_active_io_dat_actv_nz_0_67; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_68 = u_active_io_dat_actv_nz_0_68; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_69 = u_active_io_dat_actv_nz_0_69; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_70 = u_active_io_dat_actv_nz_0_70; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_71 = u_active_io_dat_actv_nz_0_71; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_72 = u_active_io_dat_actv_nz_0_72; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_73 = u_active_io_dat_actv_nz_0_73; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_74 = u_active_io_dat_actv_nz_0_74; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_75 = u_active_io_dat_actv_nz_0_75; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_76 = u_active_io_dat_actv_nz_0_76; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_77 = u_active_io_dat_actv_nz_0_77; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_78 = u_active_io_dat_actv_nz_0_78; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_79 = u_active_io_dat_actv_nz_0_79; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_80 = u_active_io_dat_actv_nz_0_80; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_81 = u_active_io_dat_actv_nz_0_81; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_82 = u_active_io_dat_actv_nz_0_82; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_83 = u_active_io_dat_actv_nz_0_83; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_84 = u_active_io_dat_actv_nz_0_84; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_85 = u_active_io_dat_actv_nz_0_85; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_86 = u_active_io_dat_actv_nz_0_86; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_87 = u_active_io_dat_actv_nz_0_87; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_88 = u_active_io_dat_actv_nz_0_88; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_89 = u_active_io_dat_actv_nz_0_89; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_90 = u_active_io_dat_actv_nz_0_90; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_91 = u_active_io_dat_actv_nz_0_91; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_92 = u_active_io_dat_actv_nz_0_92; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_93 = u_active_io_dat_actv_nz_0_93; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_94 = u_active_io_dat_actv_nz_0_94; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_95 = u_active_io_dat_actv_nz_0_95; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_96 = u_active_io_dat_actv_nz_0_96; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_97 = u_active_io_dat_actv_nz_0_97; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_98 = u_active_io_dat_actv_nz_0_98; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_99 = u_active_io_dat_actv_nz_0_99; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_100 = u_active_io_dat_actv_nz_0_100; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_101 = u_active_io_dat_actv_nz_0_101; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_102 = u_active_io_dat_actv_nz_0_102; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_103 = u_active_io_dat_actv_nz_0_103; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_104 = u_active_io_dat_actv_nz_0_104; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_105 = u_active_io_dat_actv_nz_0_105; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_106 = u_active_io_dat_actv_nz_0_106; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_107 = u_active_io_dat_actv_nz_0_107; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_108 = u_active_io_dat_actv_nz_0_108; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_109 = u_active_io_dat_actv_nz_0_109; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_110 = u_active_io_dat_actv_nz_0_110; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_111 = u_active_io_dat_actv_nz_0_111; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_112 = u_active_io_dat_actv_nz_0_112; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_113 = u_active_io_dat_actv_nz_0_113; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_114 = u_active_io_dat_actv_nz_0_114; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_115 = u_active_io_dat_actv_nz_0_115; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_116 = u_active_io_dat_actv_nz_0_116; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_117 = u_active_io_dat_actv_nz_0_117; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_118 = u_active_io_dat_actv_nz_0_118; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_119 = u_active_io_dat_actv_nz_0_119; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_120 = u_active_io_dat_actv_nz_0_120; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_121 = u_active_io_dat_actv_nz_0_121; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_122 = u_active_io_dat_actv_nz_0_122; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_123 = u_active_io_dat_actv_nz_0_123; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_124 = u_active_io_dat_actv_nz_0_124; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_125 = u_active_io_dat_actv_nz_0_125; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_126 = u_active_io_dat_actv_nz_0_126; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_nz_127 = u_active_io_dat_actv_nz_0_127; // @[NV_NVDLA_CMAC_core.scala 115:33]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_0 = u_active_io_dat_actv_pvld_0_0; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_1 = u_active_io_dat_actv_pvld_0_1; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_2 = u_active_io_dat_actv_pvld_0_2; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_3 = u_active_io_dat_actv_pvld_0_3; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_4 = u_active_io_dat_actv_pvld_0_4; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_5 = u_active_io_dat_actv_pvld_0_5; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_6 = u_active_io_dat_actv_pvld_0_6; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_7 = u_active_io_dat_actv_pvld_0_7; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_8 = u_active_io_dat_actv_pvld_0_8; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_9 = u_active_io_dat_actv_pvld_0_9; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_10 = u_active_io_dat_actv_pvld_0_10; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_11 = u_active_io_dat_actv_pvld_0_11; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_12 = u_active_io_dat_actv_pvld_0_12; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_13 = u_active_io_dat_actv_pvld_0_13; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_14 = u_active_io_dat_actv_pvld_0_14; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_15 = u_active_io_dat_actv_pvld_0_15; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_16 = u_active_io_dat_actv_pvld_0_16; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_17 = u_active_io_dat_actv_pvld_0_17; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_18 = u_active_io_dat_actv_pvld_0_18; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_19 = u_active_io_dat_actv_pvld_0_19; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_20 = u_active_io_dat_actv_pvld_0_20; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_21 = u_active_io_dat_actv_pvld_0_21; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_22 = u_active_io_dat_actv_pvld_0_22; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_23 = u_active_io_dat_actv_pvld_0_23; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_24 = u_active_io_dat_actv_pvld_0_24; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_25 = u_active_io_dat_actv_pvld_0_25; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_26 = u_active_io_dat_actv_pvld_0_26; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_27 = u_active_io_dat_actv_pvld_0_27; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_28 = u_active_io_dat_actv_pvld_0_28; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_29 = u_active_io_dat_actv_pvld_0_29; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_30 = u_active_io_dat_actv_pvld_0_30; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_31 = u_active_io_dat_actv_pvld_0_31; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_32 = u_active_io_dat_actv_pvld_0_32; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_33 = u_active_io_dat_actv_pvld_0_33; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_34 = u_active_io_dat_actv_pvld_0_34; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_35 = u_active_io_dat_actv_pvld_0_35; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_36 = u_active_io_dat_actv_pvld_0_36; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_37 = u_active_io_dat_actv_pvld_0_37; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_38 = u_active_io_dat_actv_pvld_0_38; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_39 = u_active_io_dat_actv_pvld_0_39; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_40 = u_active_io_dat_actv_pvld_0_40; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_41 = u_active_io_dat_actv_pvld_0_41; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_42 = u_active_io_dat_actv_pvld_0_42; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_43 = u_active_io_dat_actv_pvld_0_43; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_44 = u_active_io_dat_actv_pvld_0_44; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_45 = u_active_io_dat_actv_pvld_0_45; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_46 = u_active_io_dat_actv_pvld_0_46; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_47 = u_active_io_dat_actv_pvld_0_47; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_48 = u_active_io_dat_actv_pvld_0_48; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_49 = u_active_io_dat_actv_pvld_0_49; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_50 = u_active_io_dat_actv_pvld_0_50; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_51 = u_active_io_dat_actv_pvld_0_51; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_52 = u_active_io_dat_actv_pvld_0_52; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_53 = u_active_io_dat_actv_pvld_0_53; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_54 = u_active_io_dat_actv_pvld_0_54; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_55 = u_active_io_dat_actv_pvld_0_55; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_56 = u_active_io_dat_actv_pvld_0_56; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_57 = u_active_io_dat_actv_pvld_0_57; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_58 = u_active_io_dat_actv_pvld_0_58; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_59 = u_active_io_dat_actv_pvld_0_59; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_60 = u_active_io_dat_actv_pvld_0_60; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_61 = u_active_io_dat_actv_pvld_0_61; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_62 = u_active_io_dat_actv_pvld_0_62; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_63 = u_active_io_dat_actv_pvld_0_63; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_64 = u_active_io_dat_actv_pvld_0_64; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_65 = u_active_io_dat_actv_pvld_0_65; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_66 = u_active_io_dat_actv_pvld_0_66; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_67 = u_active_io_dat_actv_pvld_0_67; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_68 = u_active_io_dat_actv_pvld_0_68; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_69 = u_active_io_dat_actv_pvld_0_69; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_70 = u_active_io_dat_actv_pvld_0_70; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_71 = u_active_io_dat_actv_pvld_0_71; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_72 = u_active_io_dat_actv_pvld_0_72; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_73 = u_active_io_dat_actv_pvld_0_73; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_74 = u_active_io_dat_actv_pvld_0_74; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_75 = u_active_io_dat_actv_pvld_0_75; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_76 = u_active_io_dat_actv_pvld_0_76; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_77 = u_active_io_dat_actv_pvld_0_77; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_78 = u_active_io_dat_actv_pvld_0_78; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_79 = u_active_io_dat_actv_pvld_0_79; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_80 = u_active_io_dat_actv_pvld_0_80; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_81 = u_active_io_dat_actv_pvld_0_81; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_82 = u_active_io_dat_actv_pvld_0_82; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_83 = u_active_io_dat_actv_pvld_0_83; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_84 = u_active_io_dat_actv_pvld_0_84; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_85 = u_active_io_dat_actv_pvld_0_85; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_86 = u_active_io_dat_actv_pvld_0_86; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_87 = u_active_io_dat_actv_pvld_0_87; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_88 = u_active_io_dat_actv_pvld_0_88; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_89 = u_active_io_dat_actv_pvld_0_89; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_90 = u_active_io_dat_actv_pvld_0_90; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_91 = u_active_io_dat_actv_pvld_0_91; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_92 = u_active_io_dat_actv_pvld_0_92; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_93 = u_active_io_dat_actv_pvld_0_93; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_94 = u_active_io_dat_actv_pvld_0_94; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_95 = u_active_io_dat_actv_pvld_0_95; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_96 = u_active_io_dat_actv_pvld_0_96; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_97 = u_active_io_dat_actv_pvld_0_97; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_98 = u_active_io_dat_actv_pvld_0_98; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_99 = u_active_io_dat_actv_pvld_0_99; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_100 = u_active_io_dat_actv_pvld_0_100; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_101 = u_active_io_dat_actv_pvld_0_101; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_102 = u_active_io_dat_actv_pvld_0_102; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_103 = u_active_io_dat_actv_pvld_0_103; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_104 = u_active_io_dat_actv_pvld_0_104; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_105 = u_active_io_dat_actv_pvld_0_105; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_106 = u_active_io_dat_actv_pvld_0_106; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_107 = u_active_io_dat_actv_pvld_0_107; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_108 = u_active_io_dat_actv_pvld_0_108; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_109 = u_active_io_dat_actv_pvld_0_109; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_110 = u_active_io_dat_actv_pvld_0_110; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_111 = u_active_io_dat_actv_pvld_0_111; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_112 = u_active_io_dat_actv_pvld_0_112; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_113 = u_active_io_dat_actv_pvld_0_113; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_114 = u_active_io_dat_actv_pvld_0_114; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_115 = u_active_io_dat_actv_pvld_0_115; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_116 = u_active_io_dat_actv_pvld_0_116; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_117 = u_active_io_dat_actv_pvld_0_117; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_118 = u_active_io_dat_actv_pvld_0_118; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_119 = u_active_io_dat_actv_pvld_0_119; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_120 = u_active_io_dat_actv_pvld_0_120; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_121 = u_active_io_dat_actv_pvld_0_121; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_122 = u_active_io_dat_actv_pvld_0_122; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_123 = u_active_io_dat_actv_pvld_0_123; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_124 = u_active_io_dat_actv_pvld_0_124; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_125 = u_active_io_dat_actv_pvld_0_125; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_126 = u_active_io_dat_actv_pvld_0_126; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_dat_actv_pvld_127 = u_active_io_dat_actv_pvld_0_127; // @[NV_NVDLA_CMAC_core.scala 114:35]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_0 = u_active_io_wt_actv_data_0_0; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_1 = u_active_io_wt_actv_data_0_1; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_2 = u_active_io_wt_actv_data_0_2; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_3 = u_active_io_wt_actv_data_0_3; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_4 = u_active_io_wt_actv_data_0_4; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_5 = u_active_io_wt_actv_data_0_5; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_6 = u_active_io_wt_actv_data_0_6; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_7 = u_active_io_wt_actv_data_0_7; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_8 = u_active_io_wt_actv_data_0_8; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_9 = u_active_io_wt_actv_data_0_9; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_10 = u_active_io_wt_actv_data_0_10; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_11 = u_active_io_wt_actv_data_0_11; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_12 = u_active_io_wt_actv_data_0_12; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_13 = u_active_io_wt_actv_data_0_13; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_14 = u_active_io_wt_actv_data_0_14; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_15 = u_active_io_wt_actv_data_0_15; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_16 = u_active_io_wt_actv_data_0_16; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_17 = u_active_io_wt_actv_data_0_17; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_18 = u_active_io_wt_actv_data_0_18; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_19 = u_active_io_wt_actv_data_0_19; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_20 = u_active_io_wt_actv_data_0_20; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_21 = u_active_io_wt_actv_data_0_21; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_22 = u_active_io_wt_actv_data_0_22; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_23 = u_active_io_wt_actv_data_0_23; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_24 = u_active_io_wt_actv_data_0_24; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_25 = u_active_io_wt_actv_data_0_25; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_26 = u_active_io_wt_actv_data_0_26; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_27 = u_active_io_wt_actv_data_0_27; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_28 = u_active_io_wt_actv_data_0_28; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_29 = u_active_io_wt_actv_data_0_29; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_30 = u_active_io_wt_actv_data_0_30; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_31 = u_active_io_wt_actv_data_0_31; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_32 = u_active_io_wt_actv_data_0_32; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_33 = u_active_io_wt_actv_data_0_33; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_34 = u_active_io_wt_actv_data_0_34; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_35 = u_active_io_wt_actv_data_0_35; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_36 = u_active_io_wt_actv_data_0_36; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_37 = u_active_io_wt_actv_data_0_37; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_38 = u_active_io_wt_actv_data_0_38; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_39 = u_active_io_wt_actv_data_0_39; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_40 = u_active_io_wt_actv_data_0_40; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_41 = u_active_io_wt_actv_data_0_41; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_42 = u_active_io_wt_actv_data_0_42; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_43 = u_active_io_wt_actv_data_0_43; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_44 = u_active_io_wt_actv_data_0_44; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_45 = u_active_io_wt_actv_data_0_45; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_46 = u_active_io_wt_actv_data_0_46; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_47 = u_active_io_wt_actv_data_0_47; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_48 = u_active_io_wt_actv_data_0_48; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_49 = u_active_io_wt_actv_data_0_49; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_50 = u_active_io_wt_actv_data_0_50; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_51 = u_active_io_wt_actv_data_0_51; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_52 = u_active_io_wt_actv_data_0_52; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_53 = u_active_io_wt_actv_data_0_53; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_54 = u_active_io_wt_actv_data_0_54; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_55 = u_active_io_wt_actv_data_0_55; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_56 = u_active_io_wt_actv_data_0_56; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_57 = u_active_io_wt_actv_data_0_57; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_58 = u_active_io_wt_actv_data_0_58; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_59 = u_active_io_wt_actv_data_0_59; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_60 = u_active_io_wt_actv_data_0_60; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_61 = u_active_io_wt_actv_data_0_61; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_62 = u_active_io_wt_actv_data_0_62; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_63 = u_active_io_wt_actv_data_0_63; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_64 = u_active_io_wt_actv_data_0_64; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_65 = u_active_io_wt_actv_data_0_65; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_66 = u_active_io_wt_actv_data_0_66; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_67 = u_active_io_wt_actv_data_0_67; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_68 = u_active_io_wt_actv_data_0_68; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_69 = u_active_io_wt_actv_data_0_69; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_70 = u_active_io_wt_actv_data_0_70; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_71 = u_active_io_wt_actv_data_0_71; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_72 = u_active_io_wt_actv_data_0_72; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_73 = u_active_io_wt_actv_data_0_73; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_74 = u_active_io_wt_actv_data_0_74; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_75 = u_active_io_wt_actv_data_0_75; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_76 = u_active_io_wt_actv_data_0_76; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_77 = u_active_io_wt_actv_data_0_77; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_78 = u_active_io_wt_actv_data_0_78; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_79 = u_active_io_wt_actv_data_0_79; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_80 = u_active_io_wt_actv_data_0_80; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_81 = u_active_io_wt_actv_data_0_81; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_82 = u_active_io_wt_actv_data_0_82; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_83 = u_active_io_wt_actv_data_0_83; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_84 = u_active_io_wt_actv_data_0_84; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_85 = u_active_io_wt_actv_data_0_85; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_86 = u_active_io_wt_actv_data_0_86; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_87 = u_active_io_wt_actv_data_0_87; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_88 = u_active_io_wt_actv_data_0_88; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_89 = u_active_io_wt_actv_data_0_89; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_90 = u_active_io_wt_actv_data_0_90; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_91 = u_active_io_wt_actv_data_0_91; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_92 = u_active_io_wt_actv_data_0_92; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_93 = u_active_io_wt_actv_data_0_93; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_94 = u_active_io_wt_actv_data_0_94; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_95 = u_active_io_wt_actv_data_0_95; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_96 = u_active_io_wt_actv_data_0_96; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_97 = u_active_io_wt_actv_data_0_97; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_98 = u_active_io_wt_actv_data_0_98; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_99 = u_active_io_wt_actv_data_0_99; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_100 = u_active_io_wt_actv_data_0_100; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_101 = u_active_io_wt_actv_data_0_101; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_102 = u_active_io_wt_actv_data_0_102; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_103 = u_active_io_wt_actv_data_0_103; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_104 = u_active_io_wt_actv_data_0_104; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_105 = u_active_io_wt_actv_data_0_105; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_106 = u_active_io_wt_actv_data_0_106; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_107 = u_active_io_wt_actv_data_0_107; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_108 = u_active_io_wt_actv_data_0_108; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_109 = u_active_io_wt_actv_data_0_109; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_110 = u_active_io_wt_actv_data_0_110; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_111 = u_active_io_wt_actv_data_0_111; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_112 = u_active_io_wt_actv_data_0_112; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_113 = u_active_io_wt_actv_data_0_113; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_114 = u_active_io_wt_actv_data_0_114; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_115 = u_active_io_wt_actv_data_0_115; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_116 = u_active_io_wt_actv_data_0_116; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_117 = u_active_io_wt_actv_data_0_117; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_118 = u_active_io_wt_actv_data_0_118; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_119 = u_active_io_wt_actv_data_0_119; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_120 = u_active_io_wt_actv_data_0_120; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_121 = u_active_io_wt_actv_data_0_121; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_122 = u_active_io_wt_actv_data_0_122; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_123 = u_active_io_wt_actv_data_0_123; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_124 = u_active_io_wt_actv_data_0_124; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_125 = u_active_io_wt_actv_data_0_125; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_126 = u_active_io_wt_actv_data_0_126; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_data_127 = u_active_io_wt_actv_data_0_127; // @[NV_NVDLA_CMAC_core.scala 120:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_0 = u_active_io_wt_actv_nz_0_0; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_1 = u_active_io_wt_actv_nz_0_1; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_2 = u_active_io_wt_actv_nz_0_2; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_3 = u_active_io_wt_actv_nz_0_3; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_4 = u_active_io_wt_actv_nz_0_4; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_5 = u_active_io_wt_actv_nz_0_5; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_6 = u_active_io_wt_actv_nz_0_6; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_7 = u_active_io_wt_actv_nz_0_7; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_8 = u_active_io_wt_actv_nz_0_8; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_9 = u_active_io_wt_actv_nz_0_9; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_10 = u_active_io_wt_actv_nz_0_10; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_11 = u_active_io_wt_actv_nz_0_11; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_12 = u_active_io_wt_actv_nz_0_12; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_13 = u_active_io_wt_actv_nz_0_13; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_14 = u_active_io_wt_actv_nz_0_14; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_15 = u_active_io_wt_actv_nz_0_15; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_16 = u_active_io_wt_actv_nz_0_16; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_17 = u_active_io_wt_actv_nz_0_17; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_18 = u_active_io_wt_actv_nz_0_18; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_19 = u_active_io_wt_actv_nz_0_19; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_20 = u_active_io_wt_actv_nz_0_20; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_21 = u_active_io_wt_actv_nz_0_21; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_22 = u_active_io_wt_actv_nz_0_22; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_23 = u_active_io_wt_actv_nz_0_23; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_24 = u_active_io_wt_actv_nz_0_24; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_25 = u_active_io_wt_actv_nz_0_25; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_26 = u_active_io_wt_actv_nz_0_26; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_27 = u_active_io_wt_actv_nz_0_27; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_28 = u_active_io_wt_actv_nz_0_28; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_29 = u_active_io_wt_actv_nz_0_29; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_30 = u_active_io_wt_actv_nz_0_30; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_31 = u_active_io_wt_actv_nz_0_31; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_32 = u_active_io_wt_actv_nz_0_32; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_33 = u_active_io_wt_actv_nz_0_33; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_34 = u_active_io_wt_actv_nz_0_34; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_35 = u_active_io_wt_actv_nz_0_35; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_36 = u_active_io_wt_actv_nz_0_36; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_37 = u_active_io_wt_actv_nz_0_37; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_38 = u_active_io_wt_actv_nz_0_38; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_39 = u_active_io_wt_actv_nz_0_39; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_40 = u_active_io_wt_actv_nz_0_40; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_41 = u_active_io_wt_actv_nz_0_41; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_42 = u_active_io_wt_actv_nz_0_42; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_43 = u_active_io_wt_actv_nz_0_43; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_44 = u_active_io_wt_actv_nz_0_44; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_45 = u_active_io_wt_actv_nz_0_45; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_46 = u_active_io_wt_actv_nz_0_46; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_47 = u_active_io_wt_actv_nz_0_47; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_48 = u_active_io_wt_actv_nz_0_48; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_49 = u_active_io_wt_actv_nz_0_49; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_50 = u_active_io_wt_actv_nz_0_50; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_51 = u_active_io_wt_actv_nz_0_51; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_52 = u_active_io_wt_actv_nz_0_52; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_53 = u_active_io_wt_actv_nz_0_53; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_54 = u_active_io_wt_actv_nz_0_54; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_55 = u_active_io_wt_actv_nz_0_55; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_56 = u_active_io_wt_actv_nz_0_56; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_57 = u_active_io_wt_actv_nz_0_57; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_58 = u_active_io_wt_actv_nz_0_58; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_59 = u_active_io_wt_actv_nz_0_59; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_60 = u_active_io_wt_actv_nz_0_60; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_61 = u_active_io_wt_actv_nz_0_61; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_62 = u_active_io_wt_actv_nz_0_62; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_63 = u_active_io_wt_actv_nz_0_63; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_64 = u_active_io_wt_actv_nz_0_64; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_65 = u_active_io_wt_actv_nz_0_65; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_66 = u_active_io_wt_actv_nz_0_66; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_67 = u_active_io_wt_actv_nz_0_67; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_68 = u_active_io_wt_actv_nz_0_68; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_69 = u_active_io_wt_actv_nz_0_69; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_70 = u_active_io_wt_actv_nz_0_70; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_71 = u_active_io_wt_actv_nz_0_71; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_72 = u_active_io_wt_actv_nz_0_72; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_73 = u_active_io_wt_actv_nz_0_73; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_74 = u_active_io_wt_actv_nz_0_74; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_75 = u_active_io_wt_actv_nz_0_75; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_76 = u_active_io_wt_actv_nz_0_76; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_77 = u_active_io_wt_actv_nz_0_77; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_78 = u_active_io_wt_actv_nz_0_78; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_79 = u_active_io_wt_actv_nz_0_79; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_80 = u_active_io_wt_actv_nz_0_80; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_81 = u_active_io_wt_actv_nz_0_81; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_82 = u_active_io_wt_actv_nz_0_82; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_83 = u_active_io_wt_actv_nz_0_83; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_84 = u_active_io_wt_actv_nz_0_84; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_85 = u_active_io_wt_actv_nz_0_85; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_86 = u_active_io_wt_actv_nz_0_86; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_87 = u_active_io_wt_actv_nz_0_87; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_88 = u_active_io_wt_actv_nz_0_88; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_89 = u_active_io_wt_actv_nz_0_89; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_90 = u_active_io_wt_actv_nz_0_90; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_91 = u_active_io_wt_actv_nz_0_91; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_92 = u_active_io_wt_actv_nz_0_92; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_93 = u_active_io_wt_actv_nz_0_93; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_94 = u_active_io_wt_actv_nz_0_94; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_95 = u_active_io_wt_actv_nz_0_95; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_96 = u_active_io_wt_actv_nz_0_96; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_97 = u_active_io_wt_actv_nz_0_97; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_98 = u_active_io_wt_actv_nz_0_98; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_99 = u_active_io_wt_actv_nz_0_99; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_100 = u_active_io_wt_actv_nz_0_100; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_101 = u_active_io_wt_actv_nz_0_101; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_102 = u_active_io_wt_actv_nz_0_102; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_103 = u_active_io_wt_actv_nz_0_103; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_104 = u_active_io_wt_actv_nz_0_104; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_105 = u_active_io_wt_actv_nz_0_105; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_106 = u_active_io_wt_actv_nz_0_106; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_107 = u_active_io_wt_actv_nz_0_107; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_108 = u_active_io_wt_actv_nz_0_108; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_109 = u_active_io_wt_actv_nz_0_109; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_110 = u_active_io_wt_actv_nz_0_110; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_111 = u_active_io_wt_actv_nz_0_111; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_112 = u_active_io_wt_actv_nz_0_112; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_113 = u_active_io_wt_actv_nz_0_113; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_114 = u_active_io_wt_actv_nz_0_114; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_115 = u_active_io_wt_actv_nz_0_115; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_116 = u_active_io_wt_actv_nz_0_116; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_117 = u_active_io_wt_actv_nz_0_117; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_118 = u_active_io_wt_actv_nz_0_118; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_119 = u_active_io_wt_actv_nz_0_119; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_120 = u_active_io_wt_actv_nz_0_120; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_121 = u_active_io_wt_actv_nz_0_121; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_122 = u_active_io_wt_actv_nz_0_122; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_123 = u_active_io_wt_actv_nz_0_123; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_124 = u_active_io_wt_actv_nz_0_124; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_125 = u_active_io_wt_actv_nz_0_125; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_126 = u_active_io_wt_actv_nz_0_126; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_nz_127 = u_active_io_wt_actv_nz_0_127; // @[NV_NVDLA_CMAC_core.scala 119:32]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_0 = u_active_io_wt_actv_pvld_0_0; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_1 = u_active_io_wt_actv_pvld_0_1; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_2 = u_active_io_wt_actv_pvld_0_2; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_3 = u_active_io_wt_actv_pvld_0_3; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_4 = u_active_io_wt_actv_pvld_0_4; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_5 = u_active_io_wt_actv_pvld_0_5; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_6 = u_active_io_wt_actv_pvld_0_6; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_7 = u_active_io_wt_actv_pvld_0_7; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_8 = u_active_io_wt_actv_pvld_0_8; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_9 = u_active_io_wt_actv_pvld_0_9; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_10 = u_active_io_wt_actv_pvld_0_10; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_11 = u_active_io_wt_actv_pvld_0_11; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_12 = u_active_io_wt_actv_pvld_0_12; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_13 = u_active_io_wt_actv_pvld_0_13; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_14 = u_active_io_wt_actv_pvld_0_14; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_15 = u_active_io_wt_actv_pvld_0_15; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_16 = u_active_io_wt_actv_pvld_0_16; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_17 = u_active_io_wt_actv_pvld_0_17; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_18 = u_active_io_wt_actv_pvld_0_18; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_19 = u_active_io_wt_actv_pvld_0_19; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_20 = u_active_io_wt_actv_pvld_0_20; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_21 = u_active_io_wt_actv_pvld_0_21; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_22 = u_active_io_wt_actv_pvld_0_22; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_23 = u_active_io_wt_actv_pvld_0_23; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_24 = u_active_io_wt_actv_pvld_0_24; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_25 = u_active_io_wt_actv_pvld_0_25; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_26 = u_active_io_wt_actv_pvld_0_26; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_27 = u_active_io_wt_actv_pvld_0_27; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_28 = u_active_io_wt_actv_pvld_0_28; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_29 = u_active_io_wt_actv_pvld_0_29; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_30 = u_active_io_wt_actv_pvld_0_30; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_31 = u_active_io_wt_actv_pvld_0_31; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_32 = u_active_io_wt_actv_pvld_0_32; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_33 = u_active_io_wt_actv_pvld_0_33; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_34 = u_active_io_wt_actv_pvld_0_34; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_35 = u_active_io_wt_actv_pvld_0_35; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_36 = u_active_io_wt_actv_pvld_0_36; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_37 = u_active_io_wt_actv_pvld_0_37; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_38 = u_active_io_wt_actv_pvld_0_38; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_39 = u_active_io_wt_actv_pvld_0_39; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_40 = u_active_io_wt_actv_pvld_0_40; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_41 = u_active_io_wt_actv_pvld_0_41; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_42 = u_active_io_wt_actv_pvld_0_42; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_43 = u_active_io_wt_actv_pvld_0_43; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_44 = u_active_io_wt_actv_pvld_0_44; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_45 = u_active_io_wt_actv_pvld_0_45; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_46 = u_active_io_wt_actv_pvld_0_46; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_47 = u_active_io_wt_actv_pvld_0_47; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_48 = u_active_io_wt_actv_pvld_0_48; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_49 = u_active_io_wt_actv_pvld_0_49; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_50 = u_active_io_wt_actv_pvld_0_50; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_51 = u_active_io_wt_actv_pvld_0_51; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_52 = u_active_io_wt_actv_pvld_0_52; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_53 = u_active_io_wt_actv_pvld_0_53; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_54 = u_active_io_wt_actv_pvld_0_54; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_55 = u_active_io_wt_actv_pvld_0_55; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_56 = u_active_io_wt_actv_pvld_0_56; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_57 = u_active_io_wt_actv_pvld_0_57; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_58 = u_active_io_wt_actv_pvld_0_58; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_59 = u_active_io_wt_actv_pvld_0_59; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_60 = u_active_io_wt_actv_pvld_0_60; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_61 = u_active_io_wt_actv_pvld_0_61; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_62 = u_active_io_wt_actv_pvld_0_62; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_63 = u_active_io_wt_actv_pvld_0_63; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_64 = u_active_io_wt_actv_pvld_0_64; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_65 = u_active_io_wt_actv_pvld_0_65; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_66 = u_active_io_wt_actv_pvld_0_66; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_67 = u_active_io_wt_actv_pvld_0_67; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_68 = u_active_io_wt_actv_pvld_0_68; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_69 = u_active_io_wt_actv_pvld_0_69; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_70 = u_active_io_wt_actv_pvld_0_70; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_71 = u_active_io_wt_actv_pvld_0_71; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_72 = u_active_io_wt_actv_pvld_0_72; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_73 = u_active_io_wt_actv_pvld_0_73; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_74 = u_active_io_wt_actv_pvld_0_74; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_75 = u_active_io_wt_actv_pvld_0_75; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_76 = u_active_io_wt_actv_pvld_0_76; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_77 = u_active_io_wt_actv_pvld_0_77; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_78 = u_active_io_wt_actv_pvld_0_78; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_79 = u_active_io_wt_actv_pvld_0_79; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_80 = u_active_io_wt_actv_pvld_0_80; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_81 = u_active_io_wt_actv_pvld_0_81; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_82 = u_active_io_wt_actv_pvld_0_82; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_83 = u_active_io_wt_actv_pvld_0_83; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_84 = u_active_io_wt_actv_pvld_0_84; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_85 = u_active_io_wt_actv_pvld_0_85; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_86 = u_active_io_wt_actv_pvld_0_86; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_87 = u_active_io_wt_actv_pvld_0_87; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_88 = u_active_io_wt_actv_pvld_0_88; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_89 = u_active_io_wt_actv_pvld_0_89; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_90 = u_active_io_wt_actv_pvld_0_90; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_91 = u_active_io_wt_actv_pvld_0_91; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_92 = u_active_io_wt_actv_pvld_0_92; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_93 = u_active_io_wt_actv_pvld_0_93; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_94 = u_active_io_wt_actv_pvld_0_94; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_95 = u_active_io_wt_actv_pvld_0_95; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_96 = u_active_io_wt_actv_pvld_0_96; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_97 = u_active_io_wt_actv_pvld_0_97; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_98 = u_active_io_wt_actv_pvld_0_98; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_99 = u_active_io_wt_actv_pvld_0_99; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_100 = u_active_io_wt_actv_pvld_0_100; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_101 = u_active_io_wt_actv_pvld_0_101; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_102 = u_active_io_wt_actv_pvld_0_102; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_103 = u_active_io_wt_actv_pvld_0_103; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_104 = u_active_io_wt_actv_pvld_0_104; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_105 = u_active_io_wt_actv_pvld_0_105; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_106 = u_active_io_wt_actv_pvld_0_106; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_107 = u_active_io_wt_actv_pvld_0_107; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_108 = u_active_io_wt_actv_pvld_0_108; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_109 = u_active_io_wt_actv_pvld_0_109; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_110 = u_active_io_wt_actv_pvld_0_110; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_111 = u_active_io_wt_actv_pvld_0_111; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_112 = u_active_io_wt_actv_pvld_0_112; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_113 = u_active_io_wt_actv_pvld_0_113; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_114 = u_active_io_wt_actv_pvld_0_114; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_115 = u_active_io_wt_actv_pvld_0_115; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_116 = u_active_io_wt_actv_pvld_0_116; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_117 = u_active_io_wt_actv_pvld_0_117; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_118 = u_active_io_wt_actv_pvld_0_118; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_119 = u_active_io_wt_actv_pvld_0_119; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_120 = u_active_io_wt_actv_pvld_0_120; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_121 = u_active_io_wt_actv_pvld_0_121; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_122 = u_active_io_wt_actv_pvld_0_122; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_123 = u_active_io_wt_actv_pvld_0_123; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_124 = u_active_io_wt_actv_pvld_0_124; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_125 = u_active_io_wt_actv_pvld_0_125; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_126 = u_active_io_wt_actv_pvld_0_126; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign NV_NVDLA_CMAC_CORE_mac_io_wt_actv_pvld_127 = u_active_io_wt_actv_pvld_0_127; // @[NV_NVDLA_CMAC_core.scala 118:34]
  assign u_rt_out_clock = clock;
  assign u_rt_out_reset = reset;
  assign u_rt_out_io_out_data_0 = NV_NVDLA_CMAC_CORE_mac_io_mac_out_data; // @[NV_NVDLA_CMAC_core.scala 133:26]
  assign u_rt_out_io_out_mask_0 = NV_NVDLA_CMAC_CORE_mac_io_mac_out_pvld; // @[NV_NVDLA_CMAC_core.scala 132:26]
  assign u_rt_out_io_out_pd = out_pd; // @[NV_NVDLA_CMAC_core.scala 134:24]
  assign u_rt_out_io_out_pvld = out_pvld; // @[NV_NVDLA_CMAC_core.scala 131:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1119 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_pvld = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1122 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_pd = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_1119 <= u_rt_in_io_in_dat_pvld;
    out_pvld <= _T_1119;
    if (u_rt_in_io_in_dat_pvld) begin
      _T_1122 <= u_rt_in_io_in_dat_pd;
    end
    if (u_rt_in_io_in_dat_pvld) begin
      out_pd <= _T_1122;
    end
  end
endmodule
